module neuron64in(clk, rst, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, out);

parameter W0 = 0;
parameter W1 = 0;
parameter W2 = 0;
parameter W3 = 0;
parameter W4 = 0;
parameter W5 = 0;
parameter W6 = 0;
parameter W7 = 0;
parameter W8 = 0;
parameter W9 = 0;
parameter W10 = 0;
parameter W11 = 0;
parameter W12 = 0;
parameter W13 = 0;
parameter W14 = 0;
parameter W15 = 0;
parameter W16 = 0;
parameter W17 = 0;
parameter W18 = 0;
parameter W19 = 0;
parameter W20 = 0;
parameter W21 = 0;
parameter W22 = 0;
parameter W23 = 0;
parameter W24 = 0;
parameter W25 = 0;
parameter W26 = 0;
parameter W27 = 0;
parameter W28 = 0;
parameter W29 = 0;
parameter W30 = 0;
parameter W31 = 0;
parameter W32 = 0;
parameter W33 = 0;
parameter W34 = 0;
parameter W35 = 0;
parameter W36 = 0;
parameter W37 = 0;
parameter W38 = 0;
parameter W39 = 0;
parameter W40 = 0;
parameter W41 = 0;
parameter W42 = 0;
parameter W43 = 0;
parameter W44 = 0;
parameter W45 = 0;
parameter W46 = 0;
parameter W47 = 0;
parameter W48 = 0;
parameter W49 = 0;
parameter W50 = 0;
parameter W51 = 0;
parameter W52 = 0;
parameter W53 = 0;
parameter W54 = 0;
parameter W55 = 0;
parameter W56 = 0;
parameter W57 = 0;
parameter W58 = 0;
parameter W59 = 0;
parameter W60 = 0;
parameter W61 = 0;
parameter W62 = 0;
parameter W63 = 0;

input wire clk;
input wire rst;

input signed [15:0] in0;
input signed [15:0] in1;
input signed [15:0] in2;
input signed [15:0] in3;
input signed [15:0] in4;
input signed [15:0] in5;
input signed [15:0] in6;
input signed [15:0] in7;
input signed [15:0] in8;
input signed [15:0] in9;
input signed [15:0] in10;
input signed [15:0] in11;
input signed [15:0] in12;
input signed [15:0] in13;
input signed [15:0] in14;
input signed [15:0] in15;
input signed [15:0] in16;
input signed [15:0] in17;
input signed [15:0] in18;
input signed [15:0] in19;
input signed [15:0] in20;
input signed [15:0] in21;
input signed [15:0] in22;
input signed [15:0] in23;
input signed [15:0] in24;
input signed [15:0] in25;
input signed [15:0] in26;
input signed [15:0] in27;
input signed [15:0] in28;
input signed [15:0] in29;
input signed [15:0] in30;
input signed [15:0] in31;
input signed [15:0] in32;
input signed [15:0] in33;
input signed [15:0] in34;
input signed [15:0] in35;
input signed [15:0] in36;
input signed [15:0] in37;
input signed [15:0] in38;
input signed [15:0] in39;
input signed [15:0] in40;
input signed [15:0] in41;
input signed [15:0] in42;
input signed [15:0] in43;
input signed [15:0] in44;
input signed [15:0] in45;
input signed [15:0] in46;
input signed [15:0] in47;
input signed [15:0] in48;
input signed [15:0] in49;
input signed [15:0] in50;
input signed [15:0] in51;
input signed [15:0] in52;
input signed [15:0] in53;
input signed [15:0] in54;
input signed [15:0] in55;
input signed [15:0] in56;
input signed [15:0] in57;
input signed [15:0] in58;
input signed [15:0] in59;
input signed [15:0] in60;
input signed [15:0] in61;
input signed [15:0] in62;
input signed [15:0] in63;

output reg signed [15:0] out;

reg signed [31:0] x;
reg [31:0] abs_x;
reg [31:0] y;
always @* begin
    x = in0 * W0 / 100000 + in1 * W1 / 100000 + in2 * W2 / 100000 + in3 * W3 / 100000 + in4 * W4 / 100000 + in5 * W5 / 100000 + in6 * W6 / 100000 + in7 * W7 / 100000 + in8 * W8 / 100000 + in9 * W9 / 100000 + in10 * W10 / 100000 + in11 * W11 / 100000 + in12 * W12 / 100000 + in13 * W13 / 100000 + in14 * W14 / 100000 + in15 * W15 / 100000 + in16 * W16 / 100000 + in17 * W17 / 100000 + in18 * W18 / 100000 + in19 * W19 / 100000 + in20 * W20 / 100000 + in21 * W21 / 100000 + in22 * W22 / 100000 + in23 * W23 / 100000 + in24 * W24 / 100000 + in25 * W25 / 100000 + in26 * W26 / 100000 + in27 * W27 / 100000 + in28 * W28 / 100000 + in29 * W29 / 100000 + in30 * W30 / 100000 + in31 * W31 / 100000 + in32 * W32 / 100000 + in33 * W33 / 100000 + in34 * W34 / 100000 + in35 * W35 / 100000 + in36 * W36 / 100000 + in37 * W37 / 100000 + in38 * W38 / 100000 + in39 * W39 / 100000 + in40 * W40 / 100000 + in41 * W41 / 100000 + in42 * W42 / 100000 + in43 * W43 / 100000 + in44 * W44 / 100000 + in45 * W45 / 100000 + in46 * W46 / 100000 + in47 * W47 / 100000 + in48 * W48 / 100000 + in49 * W49 / 100000 + in50 * W50 / 100000 + in51 * W51 / 100000 + in52 * W52 / 100000 + in53 * W53 / 100000 + in54 * W54 / 100000 + in55 * W55 / 100000 + in56 * W56 / 100000 + in57 * W57 / 100000 + in58 * W58 / 100000 + in59 * W59 / 100000 + in60 * W60 / 100000 + in61 * W61 / 100000 + in62 * W62 / 100000 + in63 * W63 / 100000;
    abs_x = x < 0 ? -x : x;
    if (abs_x >= 500000) y = 100000;
    else if (abs_x >= 237500) y = 3125 * abs_x / 100000 + 84375;
    else if (abs_x >= 100000) y = 12500 * abs_x / 100000 + 62500;
    else if (abs_x >= 0) y = 25000 * abs_x / 100000 + 50000;
    out = x < 0 ? 1 - y : y;
end

endmodule

module neuron100in(clk, rst, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85, in86, in87, in88, in89, in90, in91, in92, in93, in94, in95, in96, in97, in98, in99, out);

parameter W0 = 0;
parameter W1 = 0;
parameter W2 = 0;
parameter W3 = 0;
parameter W4 = 0;
parameter W5 = 0;
parameter W6 = 0;
parameter W7 = 0;
parameter W8 = 0;
parameter W9 = 0;
parameter W10 = 0;
parameter W11 = 0;
parameter W12 = 0;
parameter W13 = 0;
parameter W14 = 0;
parameter W15 = 0;
parameter W16 = 0;
parameter W17 = 0;
parameter W18 = 0;
parameter W19 = 0;
parameter W20 = 0;
parameter W21 = 0;
parameter W22 = 0;
parameter W23 = 0;
parameter W24 = 0;
parameter W25 = 0;
parameter W26 = 0;
parameter W27 = 0;
parameter W28 = 0;
parameter W29 = 0;
parameter W30 = 0;
parameter W31 = 0;
parameter W32 = 0;
parameter W33 = 0;
parameter W34 = 0;
parameter W35 = 0;
parameter W36 = 0;
parameter W37 = 0;
parameter W38 = 0;
parameter W39 = 0;
parameter W40 = 0;
parameter W41 = 0;
parameter W42 = 0;
parameter W43 = 0;
parameter W44 = 0;
parameter W45 = 0;
parameter W46 = 0;
parameter W47 = 0;
parameter W48 = 0;
parameter W49 = 0;
parameter W50 = 0;
parameter W51 = 0;
parameter W52 = 0;
parameter W53 = 0;
parameter W54 = 0;
parameter W55 = 0;
parameter W56 = 0;
parameter W57 = 0;
parameter W58 = 0;
parameter W59 = 0;
parameter W60 = 0;
parameter W61 = 0;
parameter W62 = 0;
parameter W63 = 0;
parameter W64 = 0;
parameter W65 = 0;
parameter W66 = 0;
parameter W67 = 0;
parameter W68 = 0;
parameter W69 = 0;
parameter W70 = 0;
parameter W71 = 0;
parameter W72 = 0;
parameter W73 = 0;
parameter W74 = 0;
parameter W75 = 0;
parameter W76 = 0;
parameter W77 = 0;
parameter W78 = 0;
parameter W79 = 0;
parameter W80 = 0;
parameter W81 = 0;
parameter W82 = 0;
parameter W83 = 0;
parameter W84 = 0;
parameter W85 = 0;
parameter W86 = 0;
parameter W87 = 0;
parameter W88 = 0;
parameter W89 = 0;
parameter W90 = 0;
parameter W91 = 0;
parameter W92 = 0;
parameter W93 = 0;
parameter W94 = 0;
parameter W95 = 0;
parameter W96 = 0;
parameter W97 = 0;
parameter W98 = 0;
parameter W99 = 0;

input wire clk;
input wire rst;

input signed [15:0] in0;
input signed [15:0] in1;
input signed [15:0] in2;
input signed [15:0] in3;
input signed [15:0] in4;
input signed [15:0] in5;
input signed [15:0] in6;
input signed [15:0] in7;
input signed [15:0] in8;
input signed [15:0] in9;
input signed [15:0] in10;
input signed [15:0] in11;
input signed [15:0] in12;
input signed [15:0] in13;
input signed [15:0] in14;
input signed [15:0] in15;
input signed [15:0] in16;
input signed [15:0] in17;
input signed [15:0] in18;
input signed [15:0] in19;
input signed [15:0] in20;
input signed [15:0] in21;
input signed [15:0] in22;
input signed [15:0] in23;
input signed [15:0] in24;
input signed [15:0] in25;
input signed [15:0] in26;
input signed [15:0] in27;
input signed [15:0] in28;
input signed [15:0] in29;
input signed [15:0] in30;
input signed [15:0] in31;
input signed [15:0] in32;
input signed [15:0] in33;
input signed [15:0] in34;
input signed [15:0] in35;
input signed [15:0] in36;
input signed [15:0] in37;
input signed [15:0] in38;
input signed [15:0] in39;
input signed [15:0] in40;
input signed [15:0] in41;
input signed [15:0] in42;
input signed [15:0] in43;
input signed [15:0] in44;
input signed [15:0] in45;
input signed [15:0] in46;
input signed [15:0] in47;
input signed [15:0] in48;
input signed [15:0] in49;
input signed [15:0] in50;
input signed [15:0] in51;
input signed [15:0] in52;
input signed [15:0] in53;
input signed [15:0] in54;
input signed [15:0] in55;
input signed [15:0] in56;
input signed [15:0] in57;
input signed [15:0] in58;
input signed [15:0] in59;
input signed [15:0] in60;
input signed [15:0] in61;
input signed [15:0] in62;
input signed [15:0] in63;
input signed [15:0] in64;
input signed [15:0] in65;
input signed [15:0] in66;
input signed [15:0] in67;
input signed [15:0] in68;
input signed [15:0] in69;
input signed [15:0] in70;
input signed [15:0] in71;
input signed [15:0] in72;
input signed [15:0] in73;
input signed [15:0] in74;
input signed [15:0] in75;
input signed [15:0] in76;
input signed [15:0] in77;
input signed [15:0] in78;
input signed [15:0] in79;
input signed [15:0] in80;
input signed [15:0] in81;
input signed [15:0] in82;
input signed [15:0] in83;
input signed [15:0] in84;
input signed [15:0] in85;
input signed [15:0] in86;
input signed [15:0] in87;
input signed [15:0] in88;
input signed [15:0] in89;
input signed [15:0] in90;
input signed [15:0] in91;
input signed [15:0] in92;
input signed [15:0] in93;
input signed [15:0] in94;
input signed [15:0] in95;
input signed [15:0] in96;
input signed [15:0] in97;
input signed [15:0] in98;
input signed [15:0] in99;

output reg signed [15:0] out;

reg signed [31:0] x;
reg [31:0] abs_x;
reg [31:0] y;
always @* begin
    x = in0 * W0 / 100000 + in1 * W1 / 100000 + in2 * W2 / 100000 + in3 * W3 / 100000 + in4 * W4 / 100000 + in5 * W5 / 100000 + in6 * W6 / 100000 + in7 * W7 / 100000 + in8 * W8 / 100000 + in9 * W9 / 100000 + in10 * W10 / 100000 + in11 * W11 / 100000 + in12 * W12 / 100000 + in13 * W13 / 100000 + in14 * W14 / 100000 + in15 * W15 / 100000 + in16 * W16 / 100000 + in17 * W17 / 100000 + in18 * W18 / 100000 + in19 * W19 / 100000 + in20 * W20 / 100000 + in21 * W21 / 100000 + in22 * W22 / 100000 + in23 * W23 / 100000 + in24 * W24 / 100000 + in25 * W25 / 100000 + in26 * W26 / 100000 + in27 * W27 / 100000 + in28 * W28 / 100000 + in29 * W29 / 100000 + in30 * W30 / 100000 + in31 * W31 / 100000 + in32 * W32 / 100000 + in33 * W33 / 100000 + in34 * W34 / 100000 + in35 * W35 / 100000 + in36 * W36 / 100000 + in37 * W37 / 100000 + in38 * W38 / 100000 + in39 * W39 / 100000 + in40 * W40 / 100000 + in41 * W41 / 100000 + in42 * W42 / 100000 + in43 * W43 / 100000 + in44 * W44 / 100000 + in45 * W45 / 100000 + in46 * W46 / 100000 + in47 * W47 / 100000 + in48 * W48 / 100000 + in49 * W49 / 100000 + in50 * W50 / 100000 + in51 * W51 / 100000 + in52 * W52 / 100000 + in53 * W53 / 100000 + in54 * W54 / 100000 + in55 * W55 / 100000 + in56 * W56 / 100000 + in57 * W57 / 100000 + in58 * W58 / 100000 + in59 * W59 / 100000 + in60 * W60 / 100000 + in61 * W61 / 100000 + in62 * W62 / 100000 + in63 * W63 / 100000 + in64 * W64 / 100000 + in65 * W65 / 100000 + in66 * W66 / 100000 + in67 * W67 / 100000 + in68 * W68 / 100000 + in69 * W69 / 100000 + in70 * W70 / 100000 + in71 * W71 / 100000 + in72 * W72 / 100000 + in73 * W73 / 100000 + in74 * W74 / 100000 + in75 * W75 / 100000 + in76 * W76 / 100000 + in77 * W77 / 100000 + in78 * W78 / 100000 + in79 * W79 / 100000 + in80 * W80 / 100000 + in81 * W81 / 100000 + in82 * W82 / 100000 + in83 * W83 / 100000 + in84 * W84 / 100000 + in85 * W85 / 100000 + in86 * W86 / 100000 + in87 * W87 / 100000 + in88 * W88 / 100000 + in89 * W89 / 100000 + in90 * W90 / 100000 + in91 * W91 / 100000 + in92 * W92 / 100000 + in93 * W93 / 100000 + in94 * W94 / 100000 + in95 * W95 / 100000 + in96 * W96 / 100000 + in97 * W97 / 100000 + in98 * W98 / 100000 + in99 * W99 / 100000;
    abs_x = x < 0 ? -x : x;
    if (abs_x >= 500000) y = 100000;
    else if (abs_x >= 237500) y = 3125 * abs_x / 100000 + 84375;
    else if (abs_x >= 100000) y = 12500 * abs_x / 100000 + 62500;
    else if (abs_x >= 0) y = 25000 * abs_x / 100000 + 50000;
    out = x < 0 ? 1 - y : y;
end

endmodule

module layer64in100out(clk, rst, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, out0, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13, out14, out15, out16, out17, out18, out19, out20, out21, out22, out23, out24, out25, out26, out27, out28, out29, out30, out31, out32, out33, out34, out35, out36, out37, out38, out39, out40, out41, out42, out43, out44, out45, out46, out47, out48, out49, out50, out51, out52, out53, out54, out55, out56, out57, out58, out59, out60, out61, out62, out63, out64, out65, out66, out67, out68, out69, out70, out71, out72, out73, out74, out75, out76, out77, out78, out79, out80, out81, out82, out83, out84, out85, out86, out87, out88, out89, out90, out91, out92, out93, out94, out95, out96, out97, out98, out99);

parameter W0TO0 = 0;
parameter W0TO1 = 0;
parameter W0TO2 = 0;
parameter W0TO3 = 0;
parameter W0TO4 = 0;
parameter W0TO5 = 0;
parameter W0TO6 = 0;
parameter W0TO7 = 0;
parameter W0TO8 = 0;
parameter W0TO9 = 0;
parameter W0TO10 = 0;
parameter W0TO11 = 0;
parameter W0TO12 = 0;
parameter W0TO13 = 0;
parameter W0TO14 = 0;
parameter W0TO15 = 0;
parameter W0TO16 = 0;
parameter W0TO17 = 0;
parameter W0TO18 = 0;
parameter W0TO19 = 0;
parameter W0TO20 = 0;
parameter W0TO21 = 0;
parameter W0TO22 = 0;
parameter W0TO23 = 0;
parameter W0TO24 = 0;
parameter W0TO25 = 0;
parameter W0TO26 = 0;
parameter W0TO27 = 0;
parameter W0TO28 = 0;
parameter W0TO29 = 0;
parameter W0TO30 = 0;
parameter W0TO31 = 0;
parameter W0TO32 = 0;
parameter W0TO33 = 0;
parameter W0TO34 = 0;
parameter W0TO35 = 0;
parameter W0TO36 = 0;
parameter W0TO37 = 0;
parameter W0TO38 = 0;
parameter W0TO39 = 0;
parameter W0TO40 = 0;
parameter W0TO41 = 0;
parameter W0TO42 = 0;
parameter W0TO43 = 0;
parameter W0TO44 = 0;
parameter W0TO45 = 0;
parameter W0TO46 = 0;
parameter W0TO47 = 0;
parameter W0TO48 = 0;
parameter W0TO49 = 0;
parameter W0TO50 = 0;
parameter W0TO51 = 0;
parameter W0TO52 = 0;
parameter W0TO53 = 0;
parameter W0TO54 = 0;
parameter W0TO55 = 0;
parameter W0TO56 = 0;
parameter W0TO57 = 0;
parameter W0TO58 = 0;
parameter W0TO59 = 0;
parameter W0TO60 = 0;
parameter W0TO61 = 0;
parameter W0TO62 = 0;
parameter W0TO63 = 0;
parameter W0TO64 = 0;
parameter W0TO65 = 0;
parameter W0TO66 = 0;
parameter W0TO67 = 0;
parameter W0TO68 = 0;
parameter W0TO69 = 0;
parameter W0TO70 = 0;
parameter W0TO71 = 0;
parameter W0TO72 = 0;
parameter W0TO73 = 0;
parameter W0TO74 = 0;
parameter W0TO75 = 0;
parameter W0TO76 = 0;
parameter W0TO77 = 0;
parameter W0TO78 = 0;
parameter W0TO79 = 0;
parameter W0TO80 = 0;
parameter W0TO81 = 0;
parameter W0TO82 = 0;
parameter W0TO83 = 0;
parameter W0TO84 = 0;
parameter W0TO85 = 0;
parameter W0TO86 = 0;
parameter W0TO87 = 0;
parameter W0TO88 = 0;
parameter W0TO89 = 0;
parameter W0TO90 = 0;
parameter W0TO91 = 0;
parameter W0TO92 = 0;
parameter W0TO93 = 0;
parameter W0TO94 = 0;
parameter W0TO95 = 0;
parameter W0TO96 = 0;
parameter W0TO97 = 0;
parameter W0TO98 = 0;
parameter W0TO99 = 0;
parameter W1TO0 = 0;
parameter W1TO1 = 0;
parameter W1TO2 = 0;
parameter W1TO3 = 0;
parameter W1TO4 = 0;
parameter W1TO5 = 0;
parameter W1TO6 = 0;
parameter W1TO7 = 0;
parameter W1TO8 = 0;
parameter W1TO9 = 0;
parameter W1TO10 = 0;
parameter W1TO11 = 0;
parameter W1TO12 = 0;
parameter W1TO13 = 0;
parameter W1TO14 = 0;
parameter W1TO15 = 0;
parameter W1TO16 = 0;
parameter W1TO17 = 0;
parameter W1TO18 = 0;
parameter W1TO19 = 0;
parameter W1TO20 = 0;
parameter W1TO21 = 0;
parameter W1TO22 = 0;
parameter W1TO23 = 0;
parameter W1TO24 = 0;
parameter W1TO25 = 0;
parameter W1TO26 = 0;
parameter W1TO27 = 0;
parameter W1TO28 = 0;
parameter W1TO29 = 0;
parameter W1TO30 = 0;
parameter W1TO31 = 0;
parameter W1TO32 = 0;
parameter W1TO33 = 0;
parameter W1TO34 = 0;
parameter W1TO35 = 0;
parameter W1TO36 = 0;
parameter W1TO37 = 0;
parameter W1TO38 = 0;
parameter W1TO39 = 0;
parameter W1TO40 = 0;
parameter W1TO41 = 0;
parameter W1TO42 = 0;
parameter W1TO43 = 0;
parameter W1TO44 = 0;
parameter W1TO45 = 0;
parameter W1TO46 = 0;
parameter W1TO47 = 0;
parameter W1TO48 = 0;
parameter W1TO49 = 0;
parameter W1TO50 = 0;
parameter W1TO51 = 0;
parameter W1TO52 = 0;
parameter W1TO53 = 0;
parameter W1TO54 = 0;
parameter W1TO55 = 0;
parameter W1TO56 = 0;
parameter W1TO57 = 0;
parameter W1TO58 = 0;
parameter W1TO59 = 0;
parameter W1TO60 = 0;
parameter W1TO61 = 0;
parameter W1TO62 = 0;
parameter W1TO63 = 0;
parameter W1TO64 = 0;
parameter W1TO65 = 0;
parameter W1TO66 = 0;
parameter W1TO67 = 0;
parameter W1TO68 = 0;
parameter W1TO69 = 0;
parameter W1TO70 = 0;
parameter W1TO71 = 0;
parameter W1TO72 = 0;
parameter W1TO73 = 0;
parameter W1TO74 = 0;
parameter W1TO75 = 0;
parameter W1TO76 = 0;
parameter W1TO77 = 0;
parameter W1TO78 = 0;
parameter W1TO79 = 0;
parameter W1TO80 = 0;
parameter W1TO81 = 0;
parameter W1TO82 = 0;
parameter W1TO83 = 0;
parameter W1TO84 = 0;
parameter W1TO85 = 0;
parameter W1TO86 = 0;
parameter W1TO87 = 0;
parameter W1TO88 = 0;
parameter W1TO89 = 0;
parameter W1TO90 = 0;
parameter W1TO91 = 0;
parameter W1TO92 = 0;
parameter W1TO93 = 0;
parameter W1TO94 = 0;
parameter W1TO95 = 0;
parameter W1TO96 = 0;
parameter W1TO97 = 0;
parameter W1TO98 = 0;
parameter W1TO99 = 0;
parameter W2TO0 = 0;
parameter W2TO1 = 0;
parameter W2TO2 = 0;
parameter W2TO3 = 0;
parameter W2TO4 = 0;
parameter W2TO5 = 0;
parameter W2TO6 = 0;
parameter W2TO7 = 0;
parameter W2TO8 = 0;
parameter W2TO9 = 0;
parameter W2TO10 = 0;
parameter W2TO11 = 0;
parameter W2TO12 = 0;
parameter W2TO13 = 0;
parameter W2TO14 = 0;
parameter W2TO15 = 0;
parameter W2TO16 = 0;
parameter W2TO17 = 0;
parameter W2TO18 = 0;
parameter W2TO19 = 0;
parameter W2TO20 = 0;
parameter W2TO21 = 0;
parameter W2TO22 = 0;
parameter W2TO23 = 0;
parameter W2TO24 = 0;
parameter W2TO25 = 0;
parameter W2TO26 = 0;
parameter W2TO27 = 0;
parameter W2TO28 = 0;
parameter W2TO29 = 0;
parameter W2TO30 = 0;
parameter W2TO31 = 0;
parameter W2TO32 = 0;
parameter W2TO33 = 0;
parameter W2TO34 = 0;
parameter W2TO35 = 0;
parameter W2TO36 = 0;
parameter W2TO37 = 0;
parameter W2TO38 = 0;
parameter W2TO39 = 0;
parameter W2TO40 = 0;
parameter W2TO41 = 0;
parameter W2TO42 = 0;
parameter W2TO43 = 0;
parameter W2TO44 = 0;
parameter W2TO45 = 0;
parameter W2TO46 = 0;
parameter W2TO47 = 0;
parameter W2TO48 = 0;
parameter W2TO49 = 0;
parameter W2TO50 = 0;
parameter W2TO51 = 0;
parameter W2TO52 = 0;
parameter W2TO53 = 0;
parameter W2TO54 = 0;
parameter W2TO55 = 0;
parameter W2TO56 = 0;
parameter W2TO57 = 0;
parameter W2TO58 = 0;
parameter W2TO59 = 0;
parameter W2TO60 = 0;
parameter W2TO61 = 0;
parameter W2TO62 = 0;
parameter W2TO63 = 0;
parameter W2TO64 = 0;
parameter W2TO65 = 0;
parameter W2TO66 = 0;
parameter W2TO67 = 0;
parameter W2TO68 = 0;
parameter W2TO69 = 0;
parameter W2TO70 = 0;
parameter W2TO71 = 0;
parameter W2TO72 = 0;
parameter W2TO73 = 0;
parameter W2TO74 = 0;
parameter W2TO75 = 0;
parameter W2TO76 = 0;
parameter W2TO77 = 0;
parameter W2TO78 = 0;
parameter W2TO79 = 0;
parameter W2TO80 = 0;
parameter W2TO81 = 0;
parameter W2TO82 = 0;
parameter W2TO83 = 0;
parameter W2TO84 = 0;
parameter W2TO85 = 0;
parameter W2TO86 = 0;
parameter W2TO87 = 0;
parameter W2TO88 = 0;
parameter W2TO89 = 0;
parameter W2TO90 = 0;
parameter W2TO91 = 0;
parameter W2TO92 = 0;
parameter W2TO93 = 0;
parameter W2TO94 = 0;
parameter W2TO95 = 0;
parameter W2TO96 = 0;
parameter W2TO97 = 0;
parameter W2TO98 = 0;
parameter W2TO99 = 0;
parameter W3TO0 = 0;
parameter W3TO1 = 0;
parameter W3TO2 = 0;
parameter W3TO3 = 0;
parameter W3TO4 = 0;
parameter W3TO5 = 0;
parameter W3TO6 = 0;
parameter W3TO7 = 0;
parameter W3TO8 = 0;
parameter W3TO9 = 0;
parameter W3TO10 = 0;
parameter W3TO11 = 0;
parameter W3TO12 = 0;
parameter W3TO13 = 0;
parameter W3TO14 = 0;
parameter W3TO15 = 0;
parameter W3TO16 = 0;
parameter W3TO17 = 0;
parameter W3TO18 = 0;
parameter W3TO19 = 0;
parameter W3TO20 = 0;
parameter W3TO21 = 0;
parameter W3TO22 = 0;
parameter W3TO23 = 0;
parameter W3TO24 = 0;
parameter W3TO25 = 0;
parameter W3TO26 = 0;
parameter W3TO27 = 0;
parameter W3TO28 = 0;
parameter W3TO29 = 0;
parameter W3TO30 = 0;
parameter W3TO31 = 0;
parameter W3TO32 = 0;
parameter W3TO33 = 0;
parameter W3TO34 = 0;
parameter W3TO35 = 0;
parameter W3TO36 = 0;
parameter W3TO37 = 0;
parameter W3TO38 = 0;
parameter W3TO39 = 0;
parameter W3TO40 = 0;
parameter W3TO41 = 0;
parameter W3TO42 = 0;
parameter W3TO43 = 0;
parameter W3TO44 = 0;
parameter W3TO45 = 0;
parameter W3TO46 = 0;
parameter W3TO47 = 0;
parameter W3TO48 = 0;
parameter W3TO49 = 0;
parameter W3TO50 = 0;
parameter W3TO51 = 0;
parameter W3TO52 = 0;
parameter W3TO53 = 0;
parameter W3TO54 = 0;
parameter W3TO55 = 0;
parameter W3TO56 = 0;
parameter W3TO57 = 0;
parameter W3TO58 = 0;
parameter W3TO59 = 0;
parameter W3TO60 = 0;
parameter W3TO61 = 0;
parameter W3TO62 = 0;
parameter W3TO63 = 0;
parameter W3TO64 = 0;
parameter W3TO65 = 0;
parameter W3TO66 = 0;
parameter W3TO67 = 0;
parameter W3TO68 = 0;
parameter W3TO69 = 0;
parameter W3TO70 = 0;
parameter W3TO71 = 0;
parameter W3TO72 = 0;
parameter W3TO73 = 0;
parameter W3TO74 = 0;
parameter W3TO75 = 0;
parameter W3TO76 = 0;
parameter W3TO77 = 0;
parameter W3TO78 = 0;
parameter W3TO79 = 0;
parameter W3TO80 = 0;
parameter W3TO81 = 0;
parameter W3TO82 = 0;
parameter W3TO83 = 0;
parameter W3TO84 = 0;
parameter W3TO85 = 0;
parameter W3TO86 = 0;
parameter W3TO87 = 0;
parameter W3TO88 = 0;
parameter W3TO89 = 0;
parameter W3TO90 = 0;
parameter W3TO91 = 0;
parameter W3TO92 = 0;
parameter W3TO93 = 0;
parameter W3TO94 = 0;
parameter W3TO95 = 0;
parameter W3TO96 = 0;
parameter W3TO97 = 0;
parameter W3TO98 = 0;
parameter W3TO99 = 0;
parameter W4TO0 = 0;
parameter W4TO1 = 0;
parameter W4TO2 = 0;
parameter W4TO3 = 0;
parameter W4TO4 = 0;
parameter W4TO5 = 0;
parameter W4TO6 = 0;
parameter W4TO7 = 0;
parameter W4TO8 = 0;
parameter W4TO9 = 0;
parameter W4TO10 = 0;
parameter W4TO11 = 0;
parameter W4TO12 = 0;
parameter W4TO13 = 0;
parameter W4TO14 = 0;
parameter W4TO15 = 0;
parameter W4TO16 = 0;
parameter W4TO17 = 0;
parameter W4TO18 = 0;
parameter W4TO19 = 0;
parameter W4TO20 = 0;
parameter W4TO21 = 0;
parameter W4TO22 = 0;
parameter W4TO23 = 0;
parameter W4TO24 = 0;
parameter W4TO25 = 0;
parameter W4TO26 = 0;
parameter W4TO27 = 0;
parameter W4TO28 = 0;
parameter W4TO29 = 0;
parameter W4TO30 = 0;
parameter W4TO31 = 0;
parameter W4TO32 = 0;
parameter W4TO33 = 0;
parameter W4TO34 = 0;
parameter W4TO35 = 0;
parameter W4TO36 = 0;
parameter W4TO37 = 0;
parameter W4TO38 = 0;
parameter W4TO39 = 0;
parameter W4TO40 = 0;
parameter W4TO41 = 0;
parameter W4TO42 = 0;
parameter W4TO43 = 0;
parameter W4TO44 = 0;
parameter W4TO45 = 0;
parameter W4TO46 = 0;
parameter W4TO47 = 0;
parameter W4TO48 = 0;
parameter W4TO49 = 0;
parameter W4TO50 = 0;
parameter W4TO51 = 0;
parameter W4TO52 = 0;
parameter W4TO53 = 0;
parameter W4TO54 = 0;
parameter W4TO55 = 0;
parameter W4TO56 = 0;
parameter W4TO57 = 0;
parameter W4TO58 = 0;
parameter W4TO59 = 0;
parameter W4TO60 = 0;
parameter W4TO61 = 0;
parameter W4TO62 = 0;
parameter W4TO63 = 0;
parameter W4TO64 = 0;
parameter W4TO65 = 0;
parameter W4TO66 = 0;
parameter W4TO67 = 0;
parameter W4TO68 = 0;
parameter W4TO69 = 0;
parameter W4TO70 = 0;
parameter W4TO71 = 0;
parameter W4TO72 = 0;
parameter W4TO73 = 0;
parameter W4TO74 = 0;
parameter W4TO75 = 0;
parameter W4TO76 = 0;
parameter W4TO77 = 0;
parameter W4TO78 = 0;
parameter W4TO79 = 0;
parameter W4TO80 = 0;
parameter W4TO81 = 0;
parameter W4TO82 = 0;
parameter W4TO83 = 0;
parameter W4TO84 = 0;
parameter W4TO85 = 0;
parameter W4TO86 = 0;
parameter W4TO87 = 0;
parameter W4TO88 = 0;
parameter W4TO89 = 0;
parameter W4TO90 = 0;
parameter W4TO91 = 0;
parameter W4TO92 = 0;
parameter W4TO93 = 0;
parameter W4TO94 = 0;
parameter W4TO95 = 0;
parameter W4TO96 = 0;
parameter W4TO97 = 0;
parameter W4TO98 = 0;
parameter W4TO99 = 0;
parameter W5TO0 = 0;
parameter W5TO1 = 0;
parameter W5TO2 = 0;
parameter W5TO3 = 0;
parameter W5TO4 = 0;
parameter W5TO5 = 0;
parameter W5TO6 = 0;
parameter W5TO7 = 0;
parameter W5TO8 = 0;
parameter W5TO9 = 0;
parameter W5TO10 = 0;
parameter W5TO11 = 0;
parameter W5TO12 = 0;
parameter W5TO13 = 0;
parameter W5TO14 = 0;
parameter W5TO15 = 0;
parameter W5TO16 = 0;
parameter W5TO17 = 0;
parameter W5TO18 = 0;
parameter W5TO19 = 0;
parameter W5TO20 = 0;
parameter W5TO21 = 0;
parameter W5TO22 = 0;
parameter W5TO23 = 0;
parameter W5TO24 = 0;
parameter W5TO25 = 0;
parameter W5TO26 = 0;
parameter W5TO27 = 0;
parameter W5TO28 = 0;
parameter W5TO29 = 0;
parameter W5TO30 = 0;
parameter W5TO31 = 0;
parameter W5TO32 = 0;
parameter W5TO33 = 0;
parameter W5TO34 = 0;
parameter W5TO35 = 0;
parameter W5TO36 = 0;
parameter W5TO37 = 0;
parameter W5TO38 = 0;
parameter W5TO39 = 0;
parameter W5TO40 = 0;
parameter W5TO41 = 0;
parameter W5TO42 = 0;
parameter W5TO43 = 0;
parameter W5TO44 = 0;
parameter W5TO45 = 0;
parameter W5TO46 = 0;
parameter W5TO47 = 0;
parameter W5TO48 = 0;
parameter W5TO49 = 0;
parameter W5TO50 = 0;
parameter W5TO51 = 0;
parameter W5TO52 = 0;
parameter W5TO53 = 0;
parameter W5TO54 = 0;
parameter W5TO55 = 0;
parameter W5TO56 = 0;
parameter W5TO57 = 0;
parameter W5TO58 = 0;
parameter W5TO59 = 0;
parameter W5TO60 = 0;
parameter W5TO61 = 0;
parameter W5TO62 = 0;
parameter W5TO63 = 0;
parameter W5TO64 = 0;
parameter W5TO65 = 0;
parameter W5TO66 = 0;
parameter W5TO67 = 0;
parameter W5TO68 = 0;
parameter W5TO69 = 0;
parameter W5TO70 = 0;
parameter W5TO71 = 0;
parameter W5TO72 = 0;
parameter W5TO73 = 0;
parameter W5TO74 = 0;
parameter W5TO75 = 0;
parameter W5TO76 = 0;
parameter W5TO77 = 0;
parameter W5TO78 = 0;
parameter W5TO79 = 0;
parameter W5TO80 = 0;
parameter W5TO81 = 0;
parameter W5TO82 = 0;
parameter W5TO83 = 0;
parameter W5TO84 = 0;
parameter W5TO85 = 0;
parameter W5TO86 = 0;
parameter W5TO87 = 0;
parameter W5TO88 = 0;
parameter W5TO89 = 0;
parameter W5TO90 = 0;
parameter W5TO91 = 0;
parameter W5TO92 = 0;
parameter W5TO93 = 0;
parameter W5TO94 = 0;
parameter W5TO95 = 0;
parameter W5TO96 = 0;
parameter W5TO97 = 0;
parameter W5TO98 = 0;
parameter W5TO99 = 0;
parameter W6TO0 = 0;
parameter W6TO1 = 0;
parameter W6TO2 = 0;
parameter W6TO3 = 0;
parameter W6TO4 = 0;
parameter W6TO5 = 0;
parameter W6TO6 = 0;
parameter W6TO7 = 0;
parameter W6TO8 = 0;
parameter W6TO9 = 0;
parameter W6TO10 = 0;
parameter W6TO11 = 0;
parameter W6TO12 = 0;
parameter W6TO13 = 0;
parameter W6TO14 = 0;
parameter W6TO15 = 0;
parameter W6TO16 = 0;
parameter W6TO17 = 0;
parameter W6TO18 = 0;
parameter W6TO19 = 0;
parameter W6TO20 = 0;
parameter W6TO21 = 0;
parameter W6TO22 = 0;
parameter W6TO23 = 0;
parameter W6TO24 = 0;
parameter W6TO25 = 0;
parameter W6TO26 = 0;
parameter W6TO27 = 0;
parameter W6TO28 = 0;
parameter W6TO29 = 0;
parameter W6TO30 = 0;
parameter W6TO31 = 0;
parameter W6TO32 = 0;
parameter W6TO33 = 0;
parameter W6TO34 = 0;
parameter W6TO35 = 0;
parameter W6TO36 = 0;
parameter W6TO37 = 0;
parameter W6TO38 = 0;
parameter W6TO39 = 0;
parameter W6TO40 = 0;
parameter W6TO41 = 0;
parameter W6TO42 = 0;
parameter W6TO43 = 0;
parameter W6TO44 = 0;
parameter W6TO45 = 0;
parameter W6TO46 = 0;
parameter W6TO47 = 0;
parameter W6TO48 = 0;
parameter W6TO49 = 0;
parameter W6TO50 = 0;
parameter W6TO51 = 0;
parameter W6TO52 = 0;
parameter W6TO53 = 0;
parameter W6TO54 = 0;
parameter W6TO55 = 0;
parameter W6TO56 = 0;
parameter W6TO57 = 0;
parameter W6TO58 = 0;
parameter W6TO59 = 0;
parameter W6TO60 = 0;
parameter W6TO61 = 0;
parameter W6TO62 = 0;
parameter W6TO63 = 0;
parameter W6TO64 = 0;
parameter W6TO65 = 0;
parameter W6TO66 = 0;
parameter W6TO67 = 0;
parameter W6TO68 = 0;
parameter W6TO69 = 0;
parameter W6TO70 = 0;
parameter W6TO71 = 0;
parameter W6TO72 = 0;
parameter W6TO73 = 0;
parameter W6TO74 = 0;
parameter W6TO75 = 0;
parameter W6TO76 = 0;
parameter W6TO77 = 0;
parameter W6TO78 = 0;
parameter W6TO79 = 0;
parameter W6TO80 = 0;
parameter W6TO81 = 0;
parameter W6TO82 = 0;
parameter W6TO83 = 0;
parameter W6TO84 = 0;
parameter W6TO85 = 0;
parameter W6TO86 = 0;
parameter W6TO87 = 0;
parameter W6TO88 = 0;
parameter W6TO89 = 0;
parameter W6TO90 = 0;
parameter W6TO91 = 0;
parameter W6TO92 = 0;
parameter W6TO93 = 0;
parameter W6TO94 = 0;
parameter W6TO95 = 0;
parameter W6TO96 = 0;
parameter W6TO97 = 0;
parameter W6TO98 = 0;
parameter W6TO99 = 0;
parameter W7TO0 = 0;
parameter W7TO1 = 0;
parameter W7TO2 = 0;
parameter W7TO3 = 0;
parameter W7TO4 = 0;
parameter W7TO5 = 0;
parameter W7TO6 = 0;
parameter W7TO7 = 0;
parameter W7TO8 = 0;
parameter W7TO9 = 0;
parameter W7TO10 = 0;
parameter W7TO11 = 0;
parameter W7TO12 = 0;
parameter W7TO13 = 0;
parameter W7TO14 = 0;
parameter W7TO15 = 0;
parameter W7TO16 = 0;
parameter W7TO17 = 0;
parameter W7TO18 = 0;
parameter W7TO19 = 0;
parameter W7TO20 = 0;
parameter W7TO21 = 0;
parameter W7TO22 = 0;
parameter W7TO23 = 0;
parameter W7TO24 = 0;
parameter W7TO25 = 0;
parameter W7TO26 = 0;
parameter W7TO27 = 0;
parameter W7TO28 = 0;
parameter W7TO29 = 0;
parameter W7TO30 = 0;
parameter W7TO31 = 0;
parameter W7TO32 = 0;
parameter W7TO33 = 0;
parameter W7TO34 = 0;
parameter W7TO35 = 0;
parameter W7TO36 = 0;
parameter W7TO37 = 0;
parameter W7TO38 = 0;
parameter W7TO39 = 0;
parameter W7TO40 = 0;
parameter W7TO41 = 0;
parameter W7TO42 = 0;
parameter W7TO43 = 0;
parameter W7TO44 = 0;
parameter W7TO45 = 0;
parameter W7TO46 = 0;
parameter W7TO47 = 0;
parameter W7TO48 = 0;
parameter W7TO49 = 0;
parameter W7TO50 = 0;
parameter W7TO51 = 0;
parameter W7TO52 = 0;
parameter W7TO53 = 0;
parameter W7TO54 = 0;
parameter W7TO55 = 0;
parameter W7TO56 = 0;
parameter W7TO57 = 0;
parameter W7TO58 = 0;
parameter W7TO59 = 0;
parameter W7TO60 = 0;
parameter W7TO61 = 0;
parameter W7TO62 = 0;
parameter W7TO63 = 0;
parameter W7TO64 = 0;
parameter W7TO65 = 0;
parameter W7TO66 = 0;
parameter W7TO67 = 0;
parameter W7TO68 = 0;
parameter W7TO69 = 0;
parameter W7TO70 = 0;
parameter W7TO71 = 0;
parameter W7TO72 = 0;
parameter W7TO73 = 0;
parameter W7TO74 = 0;
parameter W7TO75 = 0;
parameter W7TO76 = 0;
parameter W7TO77 = 0;
parameter W7TO78 = 0;
parameter W7TO79 = 0;
parameter W7TO80 = 0;
parameter W7TO81 = 0;
parameter W7TO82 = 0;
parameter W7TO83 = 0;
parameter W7TO84 = 0;
parameter W7TO85 = 0;
parameter W7TO86 = 0;
parameter W7TO87 = 0;
parameter W7TO88 = 0;
parameter W7TO89 = 0;
parameter W7TO90 = 0;
parameter W7TO91 = 0;
parameter W7TO92 = 0;
parameter W7TO93 = 0;
parameter W7TO94 = 0;
parameter W7TO95 = 0;
parameter W7TO96 = 0;
parameter W7TO97 = 0;
parameter W7TO98 = 0;
parameter W7TO99 = 0;
parameter W8TO0 = 0;
parameter W8TO1 = 0;
parameter W8TO2 = 0;
parameter W8TO3 = 0;
parameter W8TO4 = 0;
parameter W8TO5 = 0;
parameter W8TO6 = 0;
parameter W8TO7 = 0;
parameter W8TO8 = 0;
parameter W8TO9 = 0;
parameter W8TO10 = 0;
parameter W8TO11 = 0;
parameter W8TO12 = 0;
parameter W8TO13 = 0;
parameter W8TO14 = 0;
parameter W8TO15 = 0;
parameter W8TO16 = 0;
parameter W8TO17 = 0;
parameter W8TO18 = 0;
parameter W8TO19 = 0;
parameter W8TO20 = 0;
parameter W8TO21 = 0;
parameter W8TO22 = 0;
parameter W8TO23 = 0;
parameter W8TO24 = 0;
parameter W8TO25 = 0;
parameter W8TO26 = 0;
parameter W8TO27 = 0;
parameter W8TO28 = 0;
parameter W8TO29 = 0;
parameter W8TO30 = 0;
parameter W8TO31 = 0;
parameter W8TO32 = 0;
parameter W8TO33 = 0;
parameter W8TO34 = 0;
parameter W8TO35 = 0;
parameter W8TO36 = 0;
parameter W8TO37 = 0;
parameter W8TO38 = 0;
parameter W8TO39 = 0;
parameter W8TO40 = 0;
parameter W8TO41 = 0;
parameter W8TO42 = 0;
parameter W8TO43 = 0;
parameter W8TO44 = 0;
parameter W8TO45 = 0;
parameter W8TO46 = 0;
parameter W8TO47 = 0;
parameter W8TO48 = 0;
parameter W8TO49 = 0;
parameter W8TO50 = 0;
parameter W8TO51 = 0;
parameter W8TO52 = 0;
parameter W8TO53 = 0;
parameter W8TO54 = 0;
parameter W8TO55 = 0;
parameter W8TO56 = 0;
parameter W8TO57 = 0;
parameter W8TO58 = 0;
parameter W8TO59 = 0;
parameter W8TO60 = 0;
parameter W8TO61 = 0;
parameter W8TO62 = 0;
parameter W8TO63 = 0;
parameter W8TO64 = 0;
parameter W8TO65 = 0;
parameter W8TO66 = 0;
parameter W8TO67 = 0;
parameter W8TO68 = 0;
parameter W8TO69 = 0;
parameter W8TO70 = 0;
parameter W8TO71 = 0;
parameter W8TO72 = 0;
parameter W8TO73 = 0;
parameter W8TO74 = 0;
parameter W8TO75 = 0;
parameter W8TO76 = 0;
parameter W8TO77 = 0;
parameter W8TO78 = 0;
parameter W8TO79 = 0;
parameter W8TO80 = 0;
parameter W8TO81 = 0;
parameter W8TO82 = 0;
parameter W8TO83 = 0;
parameter W8TO84 = 0;
parameter W8TO85 = 0;
parameter W8TO86 = 0;
parameter W8TO87 = 0;
parameter W8TO88 = 0;
parameter W8TO89 = 0;
parameter W8TO90 = 0;
parameter W8TO91 = 0;
parameter W8TO92 = 0;
parameter W8TO93 = 0;
parameter W8TO94 = 0;
parameter W8TO95 = 0;
parameter W8TO96 = 0;
parameter W8TO97 = 0;
parameter W8TO98 = 0;
parameter W8TO99 = 0;
parameter W9TO0 = 0;
parameter W9TO1 = 0;
parameter W9TO2 = 0;
parameter W9TO3 = 0;
parameter W9TO4 = 0;
parameter W9TO5 = 0;
parameter W9TO6 = 0;
parameter W9TO7 = 0;
parameter W9TO8 = 0;
parameter W9TO9 = 0;
parameter W9TO10 = 0;
parameter W9TO11 = 0;
parameter W9TO12 = 0;
parameter W9TO13 = 0;
parameter W9TO14 = 0;
parameter W9TO15 = 0;
parameter W9TO16 = 0;
parameter W9TO17 = 0;
parameter W9TO18 = 0;
parameter W9TO19 = 0;
parameter W9TO20 = 0;
parameter W9TO21 = 0;
parameter W9TO22 = 0;
parameter W9TO23 = 0;
parameter W9TO24 = 0;
parameter W9TO25 = 0;
parameter W9TO26 = 0;
parameter W9TO27 = 0;
parameter W9TO28 = 0;
parameter W9TO29 = 0;
parameter W9TO30 = 0;
parameter W9TO31 = 0;
parameter W9TO32 = 0;
parameter W9TO33 = 0;
parameter W9TO34 = 0;
parameter W9TO35 = 0;
parameter W9TO36 = 0;
parameter W9TO37 = 0;
parameter W9TO38 = 0;
parameter W9TO39 = 0;
parameter W9TO40 = 0;
parameter W9TO41 = 0;
parameter W9TO42 = 0;
parameter W9TO43 = 0;
parameter W9TO44 = 0;
parameter W9TO45 = 0;
parameter W9TO46 = 0;
parameter W9TO47 = 0;
parameter W9TO48 = 0;
parameter W9TO49 = 0;
parameter W9TO50 = 0;
parameter W9TO51 = 0;
parameter W9TO52 = 0;
parameter W9TO53 = 0;
parameter W9TO54 = 0;
parameter W9TO55 = 0;
parameter W9TO56 = 0;
parameter W9TO57 = 0;
parameter W9TO58 = 0;
parameter W9TO59 = 0;
parameter W9TO60 = 0;
parameter W9TO61 = 0;
parameter W9TO62 = 0;
parameter W9TO63 = 0;
parameter W9TO64 = 0;
parameter W9TO65 = 0;
parameter W9TO66 = 0;
parameter W9TO67 = 0;
parameter W9TO68 = 0;
parameter W9TO69 = 0;
parameter W9TO70 = 0;
parameter W9TO71 = 0;
parameter W9TO72 = 0;
parameter W9TO73 = 0;
parameter W9TO74 = 0;
parameter W9TO75 = 0;
parameter W9TO76 = 0;
parameter W9TO77 = 0;
parameter W9TO78 = 0;
parameter W9TO79 = 0;
parameter W9TO80 = 0;
parameter W9TO81 = 0;
parameter W9TO82 = 0;
parameter W9TO83 = 0;
parameter W9TO84 = 0;
parameter W9TO85 = 0;
parameter W9TO86 = 0;
parameter W9TO87 = 0;
parameter W9TO88 = 0;
parameter W9TO89 = 0;
parameter W9TO90 = 0;
parameter W9TO91 = 0;
parameter W9TO92 = 0;
parameter W9TO93 = 0;
parameter W9TO94 = 0;
parameter W9TO95 = 0;
parameter W9TO96 = 0;
parameter W9TO97 = 0;
parameter W9TO98 = 0;
parameter W9TO99 = 0;
parameter W10TO0 = 0;
parameter W10TO1 = 0;
parameter W10TO2 = 0;
parameter W10TO3 = 0;
parameter W10TO4 = 0;
parameter W10TO5 = 0;
parameter W10TO6 = 0;
parameter W10TO7 = 0;
parameter W10TO8 = 0;
parameter W10TO9 = 0;
parameter W10TO10 = 0;
parameter W10TO11 = 0;
parameter W10TO12 = 0;
parameter W10TO13 = 0;
parameter W10TO14 = 0;
parameter W10TO15 = 0;
parameter W10TO16 = 0;
parameter W10TO17 = 0;
parameter W10TO18 = 0;
parameter W10TO19 = 0;
parameter W10TO20 = 0;
parameter W10TO21 = 0;
parameter W10TO22 = 0;
parameter W10TO23 = 0;
parameter W10TO24 = 0;
parameter W10TO25 = 0;
parameter W10TO26 = 0;
parameter W10TO27 = 0;
parameter W10TO28 = 0;
parameter W10TO29 = 0;
parameter W10TO30 = 0;
parameter W10TO31 = 0;
parameter W10TO32 = 0;
parameter W10TO33 = 0;
parameter W10TO34 = 0;
parameter W10TO35 = 0;
parameter W10TO36 = 0;
parameter W10TO37 = 0;
parameter W10TO38 = 0;
parameter W10TO39 = 0;
parameter W10TO40 = 0;
parameter W10TO41 = 0;
parameter W10TO42 = 0;
parameter W10TO43 = 0;
parameter W10TO44 = 0;
parameter W10TO45 = 0;
parameter W10TO46 = 0;
parameter W10TO47 = 0;
parameter W10TO48 = 0;
parameter W10TO49 = 0;
parameter W10TO50 = 0;
parameter W10TO51 = 0;
parameter W10TO52 = 0;
parameter W10TO53 = 0;
parameter W10TO54 = 0;
parameter W10TO55 = 0;
parameter W10TO56 = 0;
parameter W10TO57 = 0;
parameter W10TO58 = 0;
parameter W10TO59 = 0;
parameter W10TO60 = 0;
parameter W10TO61 = 0;
parameter W10TO62 = 0;
parameter W10TO63 = 0;
parameter W10TO64 = 0;
parameter W10TO65 = 0;
parameter W10TO66 = 0;
parameter W10TO67 = 0;
parameter W10TO68 = 0;
parameter W10TO69 = 0;
parameter W10TO70 = 0;
parameter W10TO71 = 0;
parameter W10TO72 = 0;
parameter W10TO73 = 0;
parameter W10TO74 = 0;
parameter W10TO75 = 0;
parameter W10TO76 = 0;
parameter W10TO77 = 0;
parameter W10TO78 = 0;
parameter W10TO79 = 0;
parameter W10TO80 = 0;
parameter W10TO81 = 0;
parameter W10TO82 = 0;
parameter W10TO83 = 0;
parameter W10TO84 = 0;
parameter W10TO85 = 0;
parameter W10TO86 = 0;
parameter W10TO87 = 0;
parameter W10TO88 = 0;
parameter W10TO89 = 0;
parameter W10TO90 = 0;
parameter W10TO91 = 0;
parameter W10TO92 = 0;
parameter W10TO93 = 0;
parameter W10TO94 = 0;
parameter W10TO95 = 0;
parameter W10TO96 = 0;
parameter W10TO97 = 0;
parameter W10TO98 = 0;
parameter W10TO99 = 0;
parameter W11TO0 = 0;
parameter W11TO1 = 0;
parameter W11TO2 = 0;
parameter W11TO3 = 0;
parameter W11TO4 = 0;
parameter W11TO5 = 0;
parameter W11TO6 = 0;
parameter W11TO7 = 0;
parameter W11TO8 = 0;
parameter W11TO9 = 0;
parameter W11TO10 = 0;
parameter W11TO11 = 0;
parameter W11TO12 = 0;
parameter W11TO13 = 0;
parameter W11TO14 = 0;
parameter W11TO15 = 0;
parameter W11TO16 = 0;
parameter W11TO17 = 0;
parameter W11TO18 = 0;
parameter W11TO19 = 0;
parameter W11TO20 = 0;
parameter W11TO21 = 0;
parameter W11TO22 = 0;
parameter W11TO23 = 0;
parameter W11TO24 = 0;
parameter W11TO25 = 0;
parameter W11TO26 = 0;
parameter W11TO27 = 0;
parameter W11TO28 = 0;
parameter W11TO29 = 0;
parameter W11TO30 = 0;
parameter W11TO31 = 0;
parameter W11TO32 = 0;
parameter W11TO33 = 0;
parameter W11TO34 = 0;
parameter W11TO35 = 0;
parameter W11TO36 = 0;
parameter W11TO37 = 0;
parameter W11TO38 = 0;
parameter W11TO39 = 0;
parameter W11TO40 = 0;
parameter W11TO41 = 0;
parameter W11TO42 = 0;
parameter W11TO43 = 0;
parameter W11TO44 = 0;
parameter W11TO45 = 0;
parameter W11TO46 = 0;
parameter W11TO47 = 0;
parameter W11TO48 = 0;
parameter W11TO49 = 0;
parameter W11TO50 = 0;
parameter W11TO51 = 0;
parameter W11TO52 = 0;
parameter W11TO53 = 0;
parameter W11TO54 = 0;
parameter W11TO55 = 0;
parameter W11TO56 = 0;
parameter W11TO57 = 0;
parameter W11TO58 = 0;
parameter W11TO59 = 0;
parameter W11TO60 = 0;
parameter W11TO61 = 0;
parameter W11TO62 = 0;
parameter W11TO63 = 0;
parameter W11TO64 = 0;
parameter W11TO65 = 0;
parameter W11TO66 = 0;
parameter W11TO67 = 0;
parameter W11TO68 = 0;
parameter W11TO69 = 0;
parameter W11TO70 = 0;
parameter W11TO71 = 0;
parameter W11TO72 = 0;
parameter W11TO73 = 0;
parameter W11TO74 = 0;
parameter W11TO75 = 0;
parameter W11TO76 = 0;
parameter W11TO77 = 0;
parameter W11TO78 = 0;
parameter W11TO79 = 0;
parameter W11TO80 = 0;
parameter W11TO81 = 0;
parameter W11TO82 = 0;
parameter W11TO83 = 0;
parameter W11TO84 = 0;
parameter W11TO85 = 0;
parameter W11TO86 = 0;
parameter W11TO87 = 0;
parameter W11TO88 = 0;
parameter W11TO89 = 0;
parameter W11TO90 = 0;
parameter W11TO91 = 0;
parameter W11TO92 = 0;
parameter W11TO93 = 0;
parameter W11TO94 = 0;
parameter W11TO95 = 0;
parameter W11TO96 = 0;
parameter W11TO97 = 0;
parameter W11TO98 = 0;
parameter W11TO99 = 0;
parameter W12TO0 = 0;
parameter W12TO1 = 0;
parameter W12TO2 = 0;
parameter W12TO3 = 0;
parameter W12TO4 = 0;
parameter W12TO5 = 0;
parameter W12TO6 = 0;
parameter W12TO7 = 0;
parameter W12TO8 = 0;
parameter W12TO9 = 0;
parameter W12TO10 = 0;
parameter W12TO11 = 0;
parameter W12TO12 = 0;
parameter W12TO13 = 0;
parameter W12TO14 = 0;
parameter W12TO15 = 0;
parameter W12TO16 = 0;
parameter W12TO17 = 0;
parameter W12TO18 = 0;
parameter W12TO19 = 0;
parameter W12TO20 = 0;
parameter W12TO21 = 0;
parameter W12TO22 = 0;
parameter W12TO23 = 0;
parameter W12TO24 = 0;
parameter W12TO25 = 0;
parameter W12TO26 = 0;
parameter W12TO27 = 0;
parameter W12TO28 = 0;
parameter W12TO29 = 0;
parameter W12TO30 = 0;
parameter W12TO31 = 0;
parameter W12TO32 = 0;
parameter W12TO33 = 0;
parameter W12TO34 = 0;
parameter W12TO35 = 0;
parameter W12TO36 = 0;
parameter W12TO37 = 0;
parameter W12TO38 = 0;
parameter W12TO39 = 0;
parameter W12TO40 = 0;
parameter W12TO41 = 0;
parameter W12TO42 = 0;
parameter W12TO43 = 0;
parameter W12TO44 = 0;
parameter W12TO45 = 0;
parameter W12TO46 = 0;
parameter W12TO47 = 0;
parameter W12TO48 = 0;
parameter W12TO49 = 0;
parameter W12TO50 = 0;
parameter W12TO51 = 0;
parameter W12TO52 = 0;
parameter W12TO53 = 0;
parameter W12TO54 = 0;
parameter W12TO55 = 0;
parameter W12TO56 = 0;
parameter W12TO57 = 0;
parameter W12TO58 = 0;
parameter W12TO59 = 0;
parameter W12TO60 = 0;
parameter W12TO61 = 0;
parameter W12TO62 = 0;
parameter W12TO63 = 0;
parameter W12TO64 = 0;
parameter W12TO65 = 0;
parameter W12TO66 = 0;
parameter W12TO67 = 0;
parameter W12TO68 = 0;
parameter W12TO69 = 0;
parameter W12TO70 = 0;
parameter W12TO71 = 0;
parameter W12TO72 = 0;
parameter W12TO73 = 0;
parameter W12TO74 = 0;
parameter W12TO75 = 0;
parameter W12TO76 = 0;
parameter W12TO77 = 0;
parameter W12TO78 = 0;
parameter W12TO79 = 0;
parameter W12TO80 = 0;
parameter W12TO81 = 0;
parameter W12TO82 = 0;
parameter W12TO83 = 0;
parameter W12TO84 = 0;
parameter W12TO85 = 0;
parameter W12TO86 = 0;
parameter W12TO87 = 0;
parameter W12TO88 = 0;
parameter W12TO89 = 0;
parameter W12TO90 = 0;
parameter W12TO91 = 0;
parameter W12TO92 = 0;
parameter W12TO93 = 0;
parameter W12TO94 = 0;
parameter W12TO95 = 0;
parameter W12TO96 = 0;
parameter W12TO97 = 0;
parameter W12TO98 = 0;
parameter W12TO99 = 0;
parameter W13TO0 = 0;
parameter W13TO1 = 0;
parameter W13TO2 = 0;
parameter W13TO3 = 0;
parameter W13TO4 = 0;
parameter W13TO5 = 0;
parameter W13TO6 = 0;
parameter W13TO7 = 0;
parameter W13TO8 = 0;
parameter W13TO9 = 0;
parameter W13TO10 = 0;
parameter W13TO11 = 0;
parameter W13TO12 = 0;
parameter W13TO13 = 0;
parameter W13TO14 = 0;
parameter W13TO15 = 0;
parameter W13TO16 = 0;
parameter W13TO17 = 0;
parameter W13TO18 = 0;
parameter W13TO19 = 0;
parameter W13TO20 = 0;
parameter W13TO21 = 0;
parameter W13TO22 = 0;
parameter W13TO23 = 0;
parameter W13TO24 = 0;
parameter W13TO25 = 0;
parameter W13TO26 = 0;
parameter W13TO27 = 0;
parameter W13TO28 = 0;
parameter W13TO29 = 0;
parameter W13TO30 = 0;
parameter W13TO31 = 0;
parameter W13TO32 = 0;
parameter W13TO33 = 0;
parameter W13TO34 = 0;
parameter W13TO35 = 0;
parameter W13TO36 = 0;
parameter W13TO37 = 0;
parameter W13TO38 = 0;
parameter W13TO39 = 0;
parameter W13TO40 = 0;
parameter W13TO41 = 0;
parameter W13TO42 = 0;
parameter W13TO43 = 0;
parameter W13TO44 = 0;
parameter W13TO45 = 0;
parameter W13TO46 = 0;
parameter W13TO47 = 0;
parameter W13TO48 = 0;
parameter W13TO49 = 0;
parameter W13TO50 = 0;
parameter W13TO51 = 0;
parameter W13TO52 = 0;
parameter W13TO53 = 0;
parameter W13TO54 = 0;
parameter W13TO55 = 0;
parameter W13TO56 = 0;
parameter W13TO57 = 0;
parameter W13TO58 = 0;
parameter W13TO59 = 0;
parameter W13TO60 = 0;
parameter W13TO61 = 0;
parameter W13TO62 = 0;
parameter W13TO63 = 0;
parameter W13TO64 = 0;
parameter W13TO65 = 0;
parameter W13TO66 = 0;
parameter W13TO67 = 0;
parameter W13TO68 = 0;
parameter W13TO69 = 0;
parameter W13TO70 = 0;
parameter W13TO71 = 0;
parameter W13TO72 = 0;
parameter W13TO73 = 0;
parameter W13TO74 = 0;
parameter W13TO75 = 0;
parameter W13TO76 = 0;
parameter W13TO77 = 0;
parameter W13TO78 = 0;
parameter W13TO79 = 0;
parameter W13TO80 = 0;
parameter W13TO81 = 0;
parameter W13TO82 = 0;
parameter W13TO83 = 0;
parameter W13TO84 = 0;
parameter W13TO85 = 0;
parameter W13TO86 = 0;
parameter W13TO87 = 0;
parameter W13TO88 = 0;
parameter W13TO89 = 0;
parameter W13TO90 = 0;
parameter W13TO91 = 0;
parameter W13TO92 = 0;
parameter W13TO93 = 0;
parameter W13TO94 = 0;
parameter W13TO95 = 0;
parameter W13TO96 = 0;
parameter W13TO97 = 0;
parameter W13TO98 = 0;
parameter W13TO99 = 0;
parameter W14TO0 = 0;
parameter W14TO1 = 0;
parameter W14TO2 = 0;
parameter W14TO3 = 0;
parameter W14TO4 = 0;
parameter W14TO5 = 0;
parameter W14TO6 = 0;
parameter W14TO7 = 0;
parameter W14TO8 = 0;
parameter W14TO9 = 0;
parameter W14TO10 = 0;
parameter W14TO11 = 0;
parameter W14TO12 = 0;
parameter W14TO13 = 0;
parameter W14TO14 = 0;
parameter W14TO15 = 0;
parameter W14TO16 = 0;
parameter W14TO17 = 0;
parameter W14TO18 = 0;
parameter W14TO19 = 0;
parameter W14TO20 = 0;
parameter W14TO21 = 0;
parameter W14TO22 = 0;
parameter W14TO23 = 0;
parameter W14TO24 = 0;
parameter W14TO25 = 0;
parameter W14TO26 = 0;
parameter W14TO27 = 0;
parameter W14TO28 = 0;
parameter W14TO29 = 0;
parameter W14TO30 = 0;
parameter W14TO31 = 0;
parameter W14TO32 = 0;
parameter W14TO33 = 0;
parameter W14TO34 = 0;
parameter W14TO35 = 0;
parameter W14TO36 = 0;
parameter W14TO37 = 0;
parameter W14TO38 = 0;
parameter W14TO39 = 0;
parameter W14TO40 = 0;
parameter W14TO41 = 0;
parameter W14TO42 = 0;
parameter W14TO43 = 0;
parameter W14TO44 = 0;
parameter W14TO45 = 0;
parameter W14TO46 = 0;
parameter W14TO47 = 0;
parameter W14TO48 = 0;
parameter W14TO49 = 0;
parameter W14TO50 = 0;
parameter W14TO51 = 0;
parameter W14TO52 = 0;
parameter W14TO53 = 0;
parameter W14TO54 = 0;
parameter W14TO55 = 0;
parameter W14TO56 = 0;
parameter W14TO57 = 0;
parameter W14TO58 = 0;
parameter W14TO59 = 0;
parameter W14TO60 = 0;
parameter W14TO61 = 0;
parameter W14TO62 = 0;
parameter W14TO63 = 0;
parameter W14TO64 = 0;
parameter W14TO65 = 0;
parameter W14TO66 = 0;
parameter W14TO67 = 0;
parameter W14TO68 = 0;
parameter W14TO69 = 0;
parameter W14TO70 = 0;
parameter W14TO71 = 0;
parameter W14TO72 = 0;
parameter W14TO73 = 0;
parameter W14TO74 = 0;
parameter W14TO75 = 0;
parameter W14TO76 = 0;
parameter W14TO77 = 0;
parameter W14TO78 = 0;
parameter W14TO79 = 0;
parameter W14TO80 = 0;
parameter W14TO81 = 0;
parameter W14TO82 = 0;
parameter W14TO83 = 0;
parameter W14TO84 = 0;
parameter W14TO85 = 0;
parameter W14TO86 = 0;
parameter W14TO87 = 0;
parameter W14TO88 = 0;
parameter W14TO89 = 0;
parameter W14TO90 = 0;
parameter W14TO91 = 0;
parameter W14TO92 = 0;
parameter W14TO93 = 0;
parameter W14TO94 = 0;
parameter W14TO95 = 0;
parameter W14TO96 = 0;
parameter W14TO97 = 0;
parameter W14TO98 = 0;
parameter W14TO99 = 0;
parameter W15TO0 = 0;
parameter W15TO1 = 0;
parameter W15TO2 = 0;
parameter W15TO3 = 0;
parameter W15TO4 = 0;
parameter W15TO5 = 0;
parameter W15TO6 = 0;
parameter W15TO7 = 0;
parameter W15TO8 = 0;
parameter W15TO9 = 0;
parameter W15TO10 = 0;
parameter W15TO11 = 0;
parameter W15TO12 = 0;
parameter W15TO13 = 0;
parameter W15TO14 = 0;
parameter W15TO15 = 0;
parameter W15TO16 = 0;
parameter W15TO17 = 0;
parameter W15TO18 = 0;
parameter W15TO19 = 0;
parameter W15TO20 = 0;
parameter W15TO21 = 0;
parameter W15TO22 = 0;
parameter W15TO23 = 0;
parameter W15TO24 = 0;
parameter W15TO25 = 0;
parameter W15TO26 = 0;
parameter W15TO27 = 0;
parameter W15TO28 = 0;
parameter W15TO29 = 0;
parameter W15TO30 = 0;
parameter W15TO31 = 0;
parameter W15TO32 = 0;
parameter W15TO33 = 0;
parameter W15TO34 = 0;
parameter W15TO35 = 0;
parameter W15TO36 = 0;
parameter W15TO37 = 0;
parameter W15TO38 = 0;
parameter W15TO39 = 0;
parameter W15TO40 = 0;
parameter W15TO41 = 0;
parameter W15TO42 = 0;
parameter W15TO43 = 0;
parameter W15TO44 = 0;
parameter W15TO45 = 0;
parameter W15TO46 = 0;
parameter W15TO47 = 0;
parameter W15TO48 = 0;
parameter W15TO49 = 0;
parameter W15TO50 = 0;
parameter W15TO51 = 0;
parameter W15TO52 = 0;
parameter W15TO53 = 0;
parameter W15TO54 = 0;
parameter W15TO55 = 0;
parameter W15TO56 = 0;
parameter W15TO57 = 0;
parameter W15TO58 = 0;
parameter W15TO59 = 0;
parameter W15TO60 = 0;
parameter W15TO61 = 0;
parameter W15TO62 = 0;
parameter W15TO63 = 0;
parameter W15TO64 = 0;
parameter W15TO65 = 0;
parameter W15TO66 = 0;
parameter W15TO67 = 0;
parameter W15TO68 = 0;
parameter W15TO69 = 0;
parameter W15TO70 = 0;
parameter W15TO71 = 0;
parameter W15TO72 = 0;
parameter W15TO73 = 0;
parameter W15TO74 = 0;
parameter W15TO75 = 0;
parameter W15TO76 = 0;
parameter W15TO77 = 0;
parameter W15TO78 = 0;
parameter W15TO79 = 0;
parameter W15TO80 = 0;
parameter W15TO81 = 0;
parameter W15TO82 = 0;
parameter W15TO83 = 0;
parameter W15TO84 = 0;
parameter W15TO85 = 0;
parameter W15TO86 = 0;
parameter W15TO87 = 0;
parameter W15TO88 = 0;
parameter W15TO89 = 0;
parameter W15TO90 = 0;
parameter W15TO91 = 0;
parameter W15TO92 = 0;
parameter W15TO93 = 0;
parameter W15TO94 = 0;
parameter W15TO95 = 0;
parameter W15TO96 = 0;
parameter W15TO97 = 0;
parameter W15TO98 = 0;
parameter W15TO99 = 0;
parameter W16TO0 = 0;
parameter W16TO1 = 0;
parameter W16TO2 = 0;
parameter W16TO3 = 0;
parameter W16TO4 = 0;
parameter W16TO5 = 0;
parameter W16TO6 = 0;
parameter W16TO7 = 0;
parameter W16TO8 = 0;
parameter W16TO9 = 0;
parameter W16TO10 = 0;
parameter W16TO11 = 0;
parameter W16TO12 = 0;
parameter W16TO13 = 0;
parameter W16TO14 = 0;
parameter W16TO15 = 0;
parameter W16TO16 = 0;
parameter W16TO17 = 0;
parameter W16TO18 = 0;
parameter W16TO19 = 0;
parameter W16TO20 = 0;
parameter W16TO21 = 0;
parameter W16TO22 = 0;
parameter W16TO23 = 0;
parameter W16TO24 = 0;
parameter W16TO25 = 0;
parameter W16TO26 = 0;
parameter W16TO27 = 0;
parameter W16TO28 = 0;
parameter W16TO29 = 0;
parameter W16TO30 = 0;
parameter W16TO31 = 0;
parameter W16TO32 = 0;
parameter W16TO33 = 0;
parameter W16TO34 = 0;
parameter W16TO35 = 0;
parameter W16TO36 = 0;
parameter W16TO37 = 0;
parameter W16TO38 = 0;
parameter W16TO39 = 0;
parameter W16TO40 = 0;
parameter W16TO41 = 0;
parameter W16TO42 = 0;
parameter W16TO43 = 0;
parameter W16TO44 = 0;
parameter W16TO45 = 0;
parameter W16TO46 = 0;
parameter W16TO47 = 0;
parameter W16TO48 = 0;
parameter W16TO49 = 0;
parameter W16TO50 = 0;
parameter W16TO51 = 0;
parameter W16TO52 = 0;
parameter W16TO53 = 0;
parameter W16TO54 = 0;
parameter W16TO55 = 0;
parameter W16TO56 = 0;
parameter W16TO57 = 0;
parameter W16TO58 = 0;
parameter W16TO59 = 0;
parameter W16TO60 = 0;
parameter W16TO61 = 0;
parameter W16TO62 = 0;
parameter W16TO63 = 0;
parameter W16TO64 = 0;
parameter W16TO65 = 0;
parameter W16TO66 = 0;
parameter W16TO67 = 0;
parameter W16TO68 = 0;
parameter W16TO69 = 0;
parameter W16TO70 = 0;
parameter W16TO71 = 0;
parameter W16TO72 = 0;
parameter W16TO73 = 0;
parameter W16TO74 = 0;
parameter W16TO75 = 0;
parameter W16TO76 = 0;
parameter W16TO77 = 0;
parameter W16TO78 = 0;
parameter W16TO79 = 0;
parameter W16TO80 = 0;
parameter W16TO81 = 0;
parameter W16TO82 = 0;
parameter W16TO83 = 0;
parameter W16TO84 = 0;
parameter W16TO85 = 0;
parameter W16TO86 = 0;
parameter W16TO87 = 0;
parameter W16TO88 = 0;
parameter W16TO89 = 0;
parameter W16TO90 = 0;
parameter W16TO91 = 0;
parameter W16TO92 = 0;
parameter W16TO93 = 0;
parameter W16TO94 = 0;
parameter W16TO95 = 0;
parameter W16TO96 = 0;
parameter W16TO97 = 0;
parameter W16TO98 = 0;
parameter W16TO99 = 0;
parameter W17TO0 = 0;
parameter W17TO1 = 0;
parameter W17TO2 = 0;
parameter W17TO3 = 0;
parameter W17TO4 = 0;
parameter W17TO5 = 0;
parameter W17TO6 = 0;
parameter W17TO7 = 0;
parameter W17TO8 = 0;
parameter W17TO9 = 0;
parameter W17TO10 = 0;
parameter W17TO11 = 0;
parameter W17TO12 = 0;
parameter W17TO13 = 0;
parameter W17TO14 = 0;
parameter W17TO15 = 0;
parameter W17TO16 = 0;
parameter W17TO17 = 0;
parameter W17TO18 = 0;
parameter W17TO19 = 0;
parameter W17TO20 = 0;
parameter W17TO21 = 0;
parameter W17TO22 = 0;
parameter W17TO23 = 0;
parameter W17TO24 = 0;
parameter W17TO25 = 0;
parameter W17TO26 = 0;
parameter W17TO27 = 0;
parameter W17TO28 = 0;
parameter W17TO29 = 0;
parameter W17TO30 = 0;
parameter W17TO31 = 0;
parameter W17TO32 = 0;
parameter W17TO33 = 0;
parameter W17TO34 = 0;
parameter W17TO35 = 0;
parameter W17TO36 = 0;
parameter W17TO37 = 0;
parameter W17TO38 = 0;
parameter W17TO39 = 0;
parameter W17TO40 = 0;
parameter W17TO41 = 0;
parameter W17TO42 = 0;
parameter W17TO43 = 0;
parameter W17TO44 = 0;
parameter W17TO45 = 0;
parameter W17TO46 = 0;
parameter W17TO47 = 0;
parameter W17TO48 = 0;
parameter W17TO49 = 0;
parameter W17TO50 = 0;
parameter W17TO51 = 0;
parameter W17TO52 = 0;
parameter W17TO53 = 0;
parameter W17TO54 = 0;
parameter W17TO55 = 0;
parameter W17TO56 = 0;
parameter W17TO57 = 0;
parameter W17TO58 = 0;
parameter W17TO59 = 0;
parameter W17TO60 = 0;
parameter W17TO61 = 0;
parameter W17TO62 = 0;
parameter W17TO63 = 0;
parameter W17TO64 = 0;
parameter W17TO65 = 0;
parameter W17TO66 = 0;
parameter W17TO67 = 0;
parameter W17TO68 = 0;
parameter W17TO69 = 0;
parameter W17TO70 = 0;
parameter W17TO71 = 0;
parameter W17TO72 = 0;
parameter W17TO73 = 0;
parameter W17TO74 = 0;
parameter W17TO75 = 0;
parameter W17TO76 = 0;
parameter W17TO77 = 0;
parameter W17TO78 = 0;
parameter W17TO79 = 0;
parameter W17TO80 = 0;
parameter W17TO81 = 0;
parameter W17TO82 = 0;
parameter W17TO83 = 0;
parameter W17TO84 = 0;
parameter W17TO85 = 0;
parameter W17TO86 = 0;
parameter W17TO87 = 0;
parameter W17TO88 = 0;
parameter W17TO89 = 0;
parameter W17TO90 = 0;
parameter W17TO91 = 0;
parameter W17TO92 = 0;
parameter W17TO93 = 0;
parameter W17TO94 = 0;
parameter W17TO95 = 0;
parameter W17TO96 = 0;
parameter W17TO97 = 0;
parameter W17TO98 = 0;
parameter W17TO99 = 0;
parameter W18TO0 = 0;
parameter W18TO1 = 0;
parameter W18TO2 = 0;
parameter W18TO3 = 0;
parameter W18TO4 = 0;
parameter W18TO5 = 0;
parameter W18TO6 = 0;
parameter W18TO7 = 0;
parameter W18TO8 = 0;
parameter W18TO9 = 0;
parameter W18TO10 = 0;
parameter W18TO11 = 0;
parameter W18TO12 = 0;
parameter W18TO13 = 0;
parameter W18TO14 = 0;
parameter W18TO15 = 0;
parameter W18TO16 = 0;
parameter W18TO17 = 0;
parameter W18TO18 = 0;
parameter W18TO19 = 0;
parameter W18TO20 = 0;
parameter W18TO21 = 0;
parameter W18TO22 = 0;
parameter W18TO23 = 0;
parameter W18TO24 = 0;
parameter W18TO25 = 0;
parameter W18TO26 = 0;
parameter W18TO27 = 0;
parameter W18TO28 = 0;
parameter W18TO29 = 0;
parameter W18TO30 = 0;
parameter W18TO31 = 0;
parameter W18TO32 = 0;
parameter W18TO33 = 0;
parameter W18TO34 = 0;
parameter W18TO35 = 0;
parameter W18TO36 = 0;
parameter W18TO37 = 0;
parameter W18TO38 = 0;
parameter W18TO39 = 0;
parameter W18TO40 = 0;
parameter W18TO41 = 0;
parameter W18TO42 = 0;
parameter W18TO43 = 0;
parameter W18TO44 = 0;
parameter W18TO45 = 0;
parameter W18TO46 = 0;
parameter W18TO47 = 0;
parameter W18TO48 = 0;
parameter W18TO49 = 0;
parameter W18TO50 = 0;
parameter W18TO51 = 0;
parameter W18TO52 = 0;
parameter W18TO53 = 0;
parameter W18TO54 = 0;
parameter W18TO55 = 0;
parameter W18TO56 = 0;
parameter W18TO57 = 0;
parameter W18TO58 = 0;
parameter W18TO59 = 0;
parameter W18TO60 = 0;
parameter W18TO61 = 0;
parameter W18TO62 = 0;
parameter W18TO63 = 0;
parameter W18TO64 = 0;
parameter W18TO65 = 0;
parameter W18TO66 = 0;
parameter W18TO67 = 0;
parameter W18TO68 = 0;
parameter W18TO69 = 0;
parameter W18TO70 = 0;
parameter W18TO71 = 0;
parameter W18TO72 = 0;
parameter W18TO73 = 0;
parameter W18TO74 = 0;
parameter W18TO75 = 0;
parameter W18TO76 = 0;
parameter W18TO77 = 0;
parameter W18TO78 = 0;
parameter W18TO79 = 0;
parameter W18TO80 = 0;
parameter W18TO81 = 0;
parameter W18TO82 = 0;
parameter W18TO83 = 0;
parameter W18TO84 = 0;
parameter W18TO85 = 0;
parameter W18TO86 = 0;
parameter W18TO87 = 0;
parameter W18TO88 = 0;
parameter W18TO89 = 0;
parameter W18TO90 = 0;
parameter W18TO91 = 0;
parameter W18TO92 = 0;
parameter W18TO93 = 0;
parameter W18TO94 = 0;
parameter W18TO95 = 0;
parameter W18TO96 = 0;
parameter W18TO97 = 0;
parameter W18TO98 = 0;
parameter W18TO99 = 0;
parameter W19TO0 = 0;
parameter W19TO1 = 0;
parameter W19TO2 = 0;
parameter W19TO3 = 0;
parameter W19TO4 = 0;
parameter W19TO5 = 0;
parameter W19TO6 = 0;
parameter W19TO7 = 0;
parameter W19TO8 = 0;
parameter W19TO9 = 0;
parameter W19TO10 = 0;
parameter W19TO11 = 0;
parameter W19TO12 = 0;
parameter W19TO13 = 0;
parameter W19TO14 = 0;
parameter W19TO15 = 0;
parameter W19TO16 = 0;
parameter W19TO17 = 0;
parameter W19TO18 = 0;
parameter W19TO19 = 0;
parameter W19TO20 = 0;
parameter W19TO21 = 0;
parameter W19TO22 = 0;
parameter W19TO23 = 0;
parameter W19TO24 = 0;
parameter W19TO25 = 0;
parameter W19TO26 = 0;
parameter W19TO27 = 0;
parameter W19TO28 = 0;
parameter W19TO29 = 0;
parameter W19TO30 = 0;
parameter W19TO31 = 0;
parameter W19TO32 = 0;
parameter W19TO33 = 0;
parameter W19TO34 = 0;
parameter W19TO35 = 0;
parameter W19TO36 = 0;
parameter W19TO37 = 0;
parameter W19TO38 = 0;
parameter W19TO39 = 0;
parameter W19TO40 = 0;
parameter W19TO41 = 0;
parameter W19TO42 = 0;
parameter W19TO43 = 0;
parameter W19TO44 = 0;
parameter W19TO45 = 0;
parameter W19TO46 = 0;
parameter W19TO47 = 0;
parameter W19TO48 = 0;
parameter W19TO49 = 0;
parameter W19TO50 = 0;
parameter W19TO51 = 0;
parameter W19TO52 = 0;
parameter W19TO53 = 0;
parameter W19TO54 = 0;
parameter W19TO55 = 0;
parameter W19TO56 = 0;
parameter W19TO57 = 0;
parameter W19TO58 = 0;
parameter W19TO59 = 0;
parameter W19TO60 = 0;
parameter W19TO61 = 0;
parameter W19TO62 = 0;
parameter W19TO63 = 0;
parameter W19TO64 = 0;
parameter W19TO65 = 0;
parameter W19TO66 = 0;
parameter W19TO67 = 0;
parameter W19TO68 = 0;
parameter W19TO69 = 0;
parameter W19TO70 = 0;
parameter W19TO71 = 0;
parameter W19TO72 = 0;
parameter W19TO73 = 0;
parameter W19TO74 = 0;
parameter W19TO75 = 0;
parameter W19TO76 = 0;
parameter W19TO77 = 0;
parameter W19TO78 = 0;
parameter W19TO79 = 0;
parameter W19TO80 = 0;
parameter W19TO81 = 0;
parameter W19TO82 = 0;
parameter W19TO83 = 0;
parameter W19TO84 = 0;
parameter W19TO85 = 0;
parameter W19TO86 = 0;
parameter W19TO87 = 0;
parameter W19TO88 = 0;
parameter W19TO89 = 0;
parameter W19TO90 = 0;
parameter W19TO91 = 0;
parameter W19TO92 = 0;
parameter W19TO93 = 0;
parameter W19TO94 = 0;
parameter W19TO95 = 0;
parameter W19TO96 = 0;
parameter W19TO97 = 0;
parameter W19TO98 = 0;
parameter W19TO99 = 0;
parameter W20TO0 = 0;
parameter W20TO1 = 0;
parameter W20TO2 = 0;
parameter W20TO3 = 0;
parameter W20TO4 = 0;
parameter W20TO5 = 0;
parameter W20TO6 = 0;
parameter W20TO7 = 0;
parameter W20TO8 = 0;
parameter W20TO9 = 0;
parameter W20TO10 = 0;
parameter W20TO11 = 0;
parameter W20TO12 = 0;
parameter W20TO13 = 0;
parameter W20TO14 = 0;
parameter W20TO15 = 0;
parameter W20TO16 = 0;
parameter W20TO17 = 0;
parameter W20TO18 = 0;
parameter W20TO19 = 0;
parameter W20TO20 = 0;
parameter W20TO21 = 0;
parameter W20TO22 = 0;
parameter W20TO23 = 0;
parameter W20TO24 = 0;
parameter W20TO25 = 0;
parameter W20TO26 = 0;
parameter W20TO27 = 0;
parameter W20TO28 = 0;
parameter W20TO29 = 0;
parameter W20TO30 = 0;
parameter W20TO31 = 0;
parameter W20TO32 = 0;
parameter W20TO33 = 0;
parameter W20TO34 = 0;
parameter W20TO35 = 0;
parameter W20TO36 = 0;
parameter W20TO37 = 0;
parameter W20TO38 = 0;
parameter W20TO39 = 0;
parameter W20TO40 = 0;
parameter W20TO41 = 0;
parameter W20TO42 = 0;
parameter W20TO43 = 0;
parameter W20TO44 = 0;
parameter W20TO45 = 0;
parameter W20TO46 = 0;
parameter W20TO47 = 0;
parameter W20TO48 = 0;
parameter W20TO49 = 0;
parameter W20TO50 = 0;
parameter W20TO51 = 0;
parameter W20TO52 = 0;
parameter W20TO53 = 0;
parameter W20TO54 = 0;
parameter W20TO55 = 0;
parameter W20TO56 = 0;
parameter W20TO57 = 0;
parameter W20TO58 = 0;
parameter W20TO59 = 0;
parameter W20TO60 = 0;
parameter W20TO61 = 0;
parameter W20TO62 = 0;
parameter W20TO63 = 0;
parameter W20TO64 = 0;
parameter W20TO65 = 0;
parameter W20TO66 = 0;
parameter W20TO67 = 0;
parameter W20TO68 = 0;
parameter W20TO69 = 0;
parameter W20TO70 = 0;
parameter W20TO71 = 0;
parameter W20TO72 = 0;
parameter W20TO73 = 0;
parameter W20TO74 = 0;
parameter W20TO75 = 0;
parameter W20TO76 = 0;
parameter W20TO77 = 0;
parameter W20TO78 = 0;
parameter W20TO79 = 0;
parameter W20TO80 = 0;
parameter W20TO81 = 0;
parameter W20TO82 = 0;
parameter W20TO83 = 0;
parameter W20TO84 = 0;
parameter W20TO85 = 0;
parameter W20TO86 = 0;
parameter W20TO87 = 0;
parameter W20TO88 = 0;
parameter W20TO89 = 0;
parameter W20TO90 = 0;
parameter W20TO91 = 0;
parameter W20TO92 = 0;
parameter W20TO93 = 0;
parameter W20TO94 = 0;
parameter W20TO95 = 0;
parameter W20TO96 = 0;
parameter W20TO97 = 0;
parameter W20TO98 = 0;
parameter W20TO99 = 0;
parameter W21TO0 = 0;
parameter W21TO1 = 0;
parameter W21TO2 = 0;
parameter W21TO3 = 0;
parameter W21TO4 = 0;
parameter W21TO5 = 0;
parameter W21TO6 = 0;
parameter W21TO7 = 0;
parameter W21TO8 = 0;
parameter W21TO9 = 0;
parameter W21TO10 = 0;
parameter W21TO11 = 0;
parameter W21TO12 = 0;
parameter W21TO13 = 0;
parameter W21TO14 = 0;
parameter W21TO15 = 0;
parameter W21TO16 = 0;
parameter W21TO17 = 0;
parameter W21TO18 = 0;
parameter W21TO19 = 0;
parameter W21TO20 = 0;
parameter W21TO21 = 0;
parameter W21TO22 = 0;
parameter W21TO23 = 0;
parameter W21TO24 = 0;
parameter W21TO25 = 0;
parameter W21TO26 = 0;
parameter W21TO27 = 0;
parameter W21TO28 = 0;
parameter W21TO29 = 0;
parameter W21TO30 = 0;
parameter W21TO31 = 0;
parameter W21TO32 = 0;
parameter W21TO33 = 0;
parameter W21TO34 = 0;
parameter W21TO35 = 0;
parameter W21TO36 = 0;
parameter W21TO37 = 0;
parameter W21TO38 = 0;
parameter W21TO39 = 0;
parameter W21TO40 = 0;
parameter W21TO41 = 0;
parameter W21TO42 = 0;
parameter W21TO43 = 0;
parameter W21TO44 = 0;
parameter W21TO45 = 0;
parameter W21TO46 = 0;
parameter W21TO47 = 0;
parameter W21TO48 = 0;
parameter W21TO49 = 0;
parameter W21TO50 = 0;
parameter W21TO51 = 0;
parameter W21TO52 = 0;
parameter W21TO53 = 0;
parameter W21TO54 = 0;
parameter W21TO55 = 0;
parameter W21TO56 = 0;
parameter W21TO57 = 0;
parameter W21TO58 = 0;
parameter W21TO59 = 0;
parameter W21TO60 = 0;
parameter W21TO61 = 0;
parameter W21TO62 = 0;
parameter W21TO63 = 0;
parameter W21TO64 = 0;
parameter W21TO65 = 0;
parameter W21TO66 = 0;
parameter W21TO67 = 0;
parameter W21TO68 = 0;
parameter W21TO69 = 0;
parameter W21TO70 = 0;
parameter W21TO71 = 0;
parameter W21TO72 = 0;
parameter W21TO73 = 0;
parameter W21TO74 = 0;
parameter W21TO75 = 0;
parameter W21TO76 = 0;
parameter W21TO77 = 0;
parameter W21TO78 = 0;
parameter W21TO79 = 0;
parameter W21TO80 = 0;
parameter W21TO81 = 0;
parameter W21TO82 = 0;
parameter W21TO83 = 0;
parameter W21TO84 = 0;
parameter W21TO85 = 0;
parameter W21TO86 = 0;
parameter W21TO87 = 0;
parameter W21TO88 = 0;
parameter W21TO89 = 0;
parameter W21TO90 = 0;
parameter W21TO91 = 0;
parameter W21TO92 = 0;
parameter W21TO93 = 0;
parameter W21TO94 = 0;
parameter W21TO95 = 0;
parameter W21TO96 = 0;
parameter W21TO97 = 0;
parameter W21TO98 = 0;
parameter W21TO99 = 0;
parameter W22TO0 = 0;
parameter W22TO1 = 0;
parameter W22TO2 = 0;
parameter W22TO3 = 0;
parameter W22TO4 = 0;
parameter W22TO5 = 0;
parameter W22TO6 = 0;
parameter W22TO7 = 0;
parameter W22TO8 = 0;
parameter W22TO9 = 0;
parameter W22TO10 = 0;
parameter W22TO11 = 0;
parameter W22TO12 = 0;
parameter W22TO13 = 0;
parameter W22TO14 = 0;
parameter W22TO15 = 0;
parameter W22TO16 = 0;
parameter W22TO17 = 0;
parameter W22TO18 = 0;
parameter W22TO19 = 0;
parameter W22TO20 = 0;
parameter W22TO21 = 0;
parameter W22TO22 = 0;
parameter W22TO23 = 0;
parameter W22TO24 = 0;
parameter W22TO25 = 0;
parameter W22TO26 = 0;
parameter W22TO27 = 0;
parameter W22TO28 = 0;
parameter W22TO29 = 0;
parameter W22TO30 = 0;
parameter W22TO31 = 0;
parameter W22TO32 = 0;
parameter W22TO33 = 0;
parameter W22TO34 = 0;
parameter W22TO35 = 0;
parameter W22TO36 = 0;
parameter W22TO37 = 0;
parameter W22TO38 = 0;
parameter W22TO39 = 0;
parameter W22TO40 = 0;
parameter W22TO41 = 0;
parameter W22TO42 = 0;
parameter W22TO43 = 0;
parameter W22TO44 = 0;
parameter W22TO45 = 0;
parameter W22TO46 = 0;
parameter W22TO47 = 0;
parameter W22TO48 = 0;
parameter W22TO49 = 0;
parameter W22TO50 = 0;
parameter W22TO51 = 0;
parameter W22TO52 = 0;
parameter W22TO53 = 0;
parameter W22TO54 = 0;
parameter W22TO55 = 0;
parameter W22TO56 = 0;
parameter W22TO57 = 0;
parameter W22TO58 = 0;
parameter W22TO59 = 0;
parameter W22TO60 = 0;
parameter W22TO61 = 0;
parameter W22TO62 = 0;
parameter W22TO63 = 0;
parameter W22TO64 = 0;
parameter W22TO65 = 0;
parameter W22TO66 = 0;
parameter W22TO67 = 0;
parameter W22TO68 = 0;
parameter W22TO69 = 0;
parameter W22TO70 = 0;
parameter W22TO71 = 0;
parameter W22TO72 = 0;
parameter W22TO73 = 0;
parameter W22TO74 = 0;
parameter W22TO75 = 0;
parameter W22TO76 = 0;
parameter W22TO77 = 0;
parameter W22TO78 = 0;
parameter W22TO79 = 0;
parameter W22TO80 = 0;
parameter W22TO81 = 0;
parameter W22TO82 = 0;
parameter W22TO83 = 0;
parameter W22TO84 = 0;
parameter W22TO85 = 0;
parameter W22TO86 = 0;
parameter W22TO87 = 0;
parameter W22TO88 = 0;
parameter W22TO89 = 0;
parameter W22TO90 = 0;
parameter W22TO91 = 0;
parameter W22TO92 = 0;
parameter W22TO93 = 0;
parameter W22TO94 = 0;
parameter W22TO95 = 0;
parameter W22TO96 = 0;
parameter W22TO97 = 0;
parameter W22TO98 = 0;
parameter W22TO99 = 0;
parameter W23TO0 = 0;
parameter W23TO1 = 0;
parameter W23TO2 = 0;
parameter W23TO3 = 0;
parameter W23TO4 = 0;
parameter W23TO5 = 0;
parameter W23TO6 = 0;
parameter W23TO7 = 0;
parameter W23TO8 = 0;
parameter W23TO9 = 0;
parameter W23TO10 = 0;
parameter W23TO11 = 0;
parameter W23TO12 = 0;
parameter W23TO13 = 0;
parameter W23TO14 = 0;
parameter W23TO15 = 0;
parameter W23TO16 = 0;
parameter W23TO17 = 0;
parameter W23TO18 = 0;
parameter W23TO19 = 0;
parameter W23TO20 = 0;
parameter W23TO21 = 0;
parameter W23TO22 = 0;
parameter W23TO23 = 0;
parameter W23TO24 = 0;
parameter W23TO25 = 0;
parameter W23TO26 = 0;
parameter W23TO27 = 0;
parameter W23TO28 = 0;
parameter W23TO29 = 0;
parameter W23TO30 = 0;
parameter W23TO31 = 0;
parameter W23TO32 = 0;
parameter W23TO33 = 0;
parameter W23TO34 = 0;
parameter W23TO35 = 0;
parameter W23TO36 = 0;
parameter W23TO37 = 0;
parameter W23TO38 = 0;
parameter W23TO39 = 0;
parameter W23TO40 = 0;
parameter W23TO41 = 0;
parameter W23TO42 = 0;
parameter W23TO43 = 0;
parameter W23TO44 = 0;
parameter W23TO45 = 0;
parameter W23TO46 = 0;
parameter W23TO47 = 0;
parameter W23TO48 = 0;
parameter W23TO49 = 0;
parameter W23TO50 = 0;
parameter W23TO51 = 0;
parameter W23TO52 = 0;
parameter W23TO53 = 0;
parameter W23TO54 = 0;
parameter W23TO55 = 0;
parameter W23TO56 = 0;
parameter W23TO57 = 0;
parameter W23TO58 = 0;
parameter W23TO59 = 0;
parameter W23TO60 = 0;
parameter W23TO61 = 0;
parameter W23TO62 = 0;
parameter W23TO63 = 0;
parameter W23TO64 = 0;
parameter W23TO65 = 0;
parameter W23TO66 = 0;
parameter W23TO67 = 0;
parameter W23TO68 = 0;
parameter W23TO69 = 0;
parameter W23TO70 = 0;
parameter W23TO71 = 0;
parameter W23TO72 = 0;
parameter W23TO73 = 0;
parameter W23TO74 = 0;
parameter W23TO75 = 0;
parameter W23TO76 = 0;
parameter W23TO77 = 0;
parameter W23TO78 = 0;
parameter W23TO79 = 0;
parameter W23TO80 = 0;
parameter W23TO81 = 0;
parameter W23TO82 = 0;
parameter W23TO83 = 0;
parameter W23TO84 = 0;
parameter W23TO85 = 0;
parameter W23TO86 = 0;
parameter W23TO87 = 0;
parameter W23TO88 = 0;
parameter W23TO89 = 0;
parameter W23TO90 = 0;
parameter W23TO91 = 0;
parameter W23TO92 = 0;
parameter W23TO93 = 0;
parameter W23TO94 = 0;
parameter W23TO95 = 0;
parameter W23TO96 = 0;
parameter W23TO97 = 0;
parameter W23TO98 = 0;
parameter W23TO99 = 0;
parameter W24TO0 = 0;
parameter W24TO1 = 0;
parameter W24TO2 = 0;
parameter W24TO3 = 0;
parameter W24TO4 = 0;
parameter W24TO5 = 0;
parameter W24TO6 = 0;
parameter W24TO7 = 0;
parameter W24TO8 = 0;
parameter W24TO9 = 0;
parameter W24TO10 = 0;
parameter W24TO11 = 0;
parameter W24TO12 = 0;
parameter W24TO13 = 0;
parameter W24TO14 = 0;
parameter W24TO15 = 0;
parameter W24TO16 = 0;
parameter W24TO17 = 0;
parameter W24TO18 = 0;
parameter W24TO19 = 0;
parameter W24TO20 = 0;
parameter W24TO21 = 0;
parameter W24TO22 = 0;
parameter W24TO23 = 0;
parameter W24TO24 = 0;
parameter W24TO25 = 0;
parameter W24TO26 = 0;
parameter W24TO27 = 0;
parameter W24TO28 = 0;
parameter W24TO29 = 0;
parameter W24TO30 = 0;
parameter W24TO31 = 0;
parameter W24TO32 = 0;
parameter W24TO33 = 0;
parameter W24TO34 = 0;
parameter W24TO35 = 0;
parameter W24TO36 = 0;
parameter W24TO37 = 0;
parameter W24TO38 = 0;
parameter W24TO39 = 0;
parameter W24TO40 = 0;
parameter W24TO41 = 0;
parameter W24TO42 = 0;
parameter W24TO43 = 0;
parameter W24TO44 = 0;
parameter W24TO45 = 0;
parameter W24TO46 = 0;
parameter W24TO47 = 0;
parameter W24TO48 = 0;
parameter W24TO49 = 0;
parameter W24TO50 = 0;
parameter W24TO51 = 0;
parameter W24TO52 = 0;
parameter W24TO53 = 0;
parameter W24TO54 = 0;
parameter W24TO55 = 0;
parameter W24TO56 = 0;
parameter W24TO57 = 0;
parameter W24TO58 = 0;
parameter W24TO59 = 0;
parameter W24TO60 = 0;
parameter W24TO61 = 0;
parameter W24TO62 = 0;
parameter W24TO63 = 0;
parameter W24TO64 = 0;
parameter W24TO65 = 0;
parameter W24TO66 = 0;
parameter W24TO67 = 0;
parameter W24TO68 = 0;
parameter W24TO69 = 0;
parameter W24TO70 = 0;
parameter W24TO71 = 0;
parameter W24TO72 = 0;
parameter W24TO73 = 0;
parameter W24TO74 = 0;
parameter W24TO75 = 0;
parameter W24TO76 = 0;
parameter W24TO77 = 0;
parameter W24TO78 = 0;
parameter W24TO79 = 0;
parameter W24TO80 = 0;
parameter W24TO81 = 0;
parameter W24TO82 = 0;
parameter W24TO83 = 0;
parameter W24TO84 = 0;
parameter W24TO85 = 0;
parameter W24TO86 = 0;
parameter W24TO87 = 0;
parameter W24TO88 = 0;
parameter W24TO89 = 0;
parameter W24TO90 = 0;
parameter W24TO91 = 0;
parameter W24TO92 = 0;
parameter W24TO93 = 0;
parameter W24TO94 = 0;
parameter W24TO95 = 0;
parameter W24TO96 = 0;
parameter W24TO97 = 0;
parameter W24TO98 = 0;
parameter W24TO99 = 0;
parameter W25TO0 = 0;
parameter W25TO1 = 0;
parameter W25TO2 = 0;
parameter W25TO3 = 0;
parameter W25TO4 = 0;
parameter W25TO5 = 0;
parameter W25TO6 = 0;
parameter W25TO7 = 0;
parameter W25TO8 = 0;
parameter W25TO9 = 0;
parameter W25TO10 = 0;
parameter W25TO11 = 0;
parameter W25TO12 = 0;
parameter W25TO13 = 0;
parameter W25TO14 = 0;
parameter W25TO15 = 0;
parameter W25TO16 = 0;
parameter W25TO17 = 0;
parameter W25TO18 = 0;
parameter W25TO19 = 0;
parameter W25TO20 = 0;
parameter W25TO21 = 0;
parameter W25TO22 = 0;
parameter W25TO23 = 0;
parameter W25TO24 = 0;
parameter W25TO25 = 0;
parameter W25TO26 = 0;
parameter W25TO27 = 0;
parameter W25TO28 = 0;
parameter W25TO29 = 0;
parameter W25TO30 = 0;
parameter W25TO31 = 0;
parameter W25TO32 = 0;
parameter W25TO33 = 0;
parameter W25TO34 = 0;
parameter W25TO35 = 0;
parameter W25TO36 = 0;
parameter W25TO37 = 0;
parameter W25TO38 = 0;
parameter W25TO39 = 0;
parameter W25TO40 = 0;
parameter W25TO41 = 0;
parameter W25TO42 = 0;
parameter W25TO43 = 0;
parameter W25TO44 = 0;
parameter W25TO45 = 0;
parameter W25TO46 = 0;
parameter W25TO47 = 0;
parameter W25TO48 = 0;
parameter W25TO49 = 0;
parameter W25TO50 = 0;
parameter W25TO51 = 0;
parameter W25TO52 = 0;
parameter W25TO53 = 0;
parameter W25TO54 = 0;
parameter W25TO55 = 0;
parameter W25TO56 = 0;
parameter W25TO57 = 0;
parameter W25TO58 = 0;
parameter W25TO59 = 0;
parameter W25TO60 = 0;
parameter W25TO61 = 0;
parameter W25TO62 = 0;
parameter W25TO63 = 0;
parameter W25TO64 = 0;
parameter W25TO65 = 0;
parameter W25TO66 = 0;
parameter W25TO67 = 0;
parameter W25TO68 = 0;
parameter W25TO69 = 0;
parameter W25TO70 = 0;
parameter W25TO71 = 0;
parameter W25TO72 = 0;
parameter W25TO73 = 0;
parameter W25TO74 = 0;
parameter W25TO75 = 0;
parameter W25TO76 = 0;
parameter W25TO77 = 0;
parameter W25TO78 = 0;
parameter W25TO79 = 0;
parameter W25TO80 = 0;
parameter W25TO81 = 0;
parameter W25TO82 = 0;
parameter W25TO83 = 0;
parameter W25TO84 = 0;
parameter W25TO85 = 0;
parameter W25TO86 = 0;
parameter W25TO87 = 0;
parameter W25TO88 = 0;
parameter W25TO89 = 0;
parameter W25TO90 = 0;
parameter W25TO91 = 0;
parameter W25TO92 = 0;
parameter W25TO93 = 0;
parameter W25TO94 = 0;
parameter W25TO95 = 0;
parameter W25TO96 = 0;
parameter W25TO97 = 0;
parameter W25TO98 = 0;
parameter W25TO99 = 0;
parameter W26TO0 = 0;
parameter W26TO1 = 0;
parameter W26TO2 = 0;
parameter W26TO3 = 0;
parameter W26TO4 = 0;
parameter W26TO5 = 0;
parameter W26TO6 = 0;
parameter W26TO7 = 0;
parameter W26TO8 = 0;
parameter W26TO9 = 0;
parameter W26TO10 = 0;
parameter W26TO11 = 0;
parameter W26TO12 = 0;
parameter W26TO13 = 0;
parameter W26TO14 = 0;
parameter W26TO15 = 0;
parameter W26TO16 = 0;
parameter W26TO17 = 0;
parameter W26TO18 = 0;
parameter W26TO19 = 0;
parameter W26TO20 = 0;
parameter W26TO21 = 0;
parameter W26TO22 = 0;
parameter W26TO23 = 0;
parameter W26TO24 = 0;
parameter W26TO25 = 0;
parameter W26TO26 = 0;
parameter W26TO27 = 0;
parameter W26TO28 = 0;
parameter W26TO29 = 0;
parameter W26TO30 = 0;
parameter W26TO31 = 0;
parameter W26TO32 = 0;
parameter W26TO33 = 0;
parameter W26TO34 = 0;
parameter W26TO35 = 0;
parameter W26TO36 = 0;
parameter W26TO37 = 0;
parameter W26TO38 = 0;
parameter W26TO39 = 0;
parameter W26TO40 = 0;
parameter W26TO41 = 0;
parameter W26TO42 = 0;
parameter W26TO43 = 0;
parameter W26TO44 = 0;
parameter W26TO45 = 0;
parameter W26TO46 = 0;
parameter W26TO47 = 0;
parameter W26TO48 = 0;
parameter W26TO49 = 0;
parameter W26TO50 = 0;
parameter W26TO51 = 0;
parameter W26TO52 = 0;
parameter W26TO53 = 0;
parameter W26TO54 = 0;
parameter W26TO55 = 0;
parameter W26TO56 = 0;
parameter W26TO57 = 0;
parameter W26TO58 = 0;
parameter W26TO59 = 0;
parameter W26TO60 = 0;
parameter W26TO61 = 0;
parameter W26TO62 = 0;
parameter W26TO63 = 0;
parameter W26TO64 = 0;
parameter W26TO65 = 0;
parameter W26TO66 = 0;
parameter W26TO67 = 0;
parameter W26TO68 = 0;
parameter W26TO69 = 0;
parameter W26TO70 = 0;
parameter W26TO71 = 0;
parameter W26TO72 = 0;
parameter W26TO73 = 0;
parameter W26TO74 = 0;
parameter W26TO75 = 0;
parameter W26TO76 = 0;
parameter W26TO77 = 0;
parameter W26TO78 = 0;
parameter W26TO79 = 0;
parameter W26TO80 = 0;
parameter W26TO81 = 0;
parameter W26TO82 = 0;
parameter W26TO83 = 0;
parameter W26TO84 = 0;
parameter W26TO85 = 0;
parameter W26TO86 = 0;
parameter W26TO87 = 0;
parameter W26TO88 = 0;
parameter W26TO89 = 0;
parameter W26TO90 = 0;
parameter W26TO91 = 0;
parameter W26TO92 = 0;
parameter W26TO93 = 0;
parameter W26TO94 = 0;
parameter W26TO95 = 0;
parameter W26TO96 = 0;
parameter W26TO97 = 0;
parameter W26TO98 = 0;
parameter W26TO99 = 0;
parameter W27TO0 = 0;
parameter W27TO1 = 0;
parameter W27TO2 = 0;
parameter W27TO3 = 0;
parameter W27TO4 = 0;
parameter W27TO5 = 0;
parameter W27TO6 = 0;
parameter W27TO7 = 0;
parameter W27TO8 = 0;
parameter W27TO9 = 0;
parameter W27TO10 = 0;
parameter W27TO11 = 0;
parameter W27TO12 = 0;
parameter W27TO13 = 0;
parameter W27TO14 = 0;
parameter W27TO15 = 0;
parameter W27TO16 = 0;
parameter W27TO17 = 0;
parameter W27TO18 = 0;
parameter W27TO19 = 0;
parameter W27TO20 = 0;
parameter W27TO21 = 0;
parameter W27TO22 = 0;
parameter W27TO23 = 0;
parameter W27TO24 = 0;
parameter W27TO25 = 0;
parameter W27TO26 = 0;
parameter W27TO27 = 0;
parameter W27TO28 = 0;
parameter W27TO29 = 0;
parameter W27TO30 = 0;
parameter W27TO31 = 0;
parameter W27TO32 = 0;
parameter W27TO33 = 0;
parameter W27TO34 = 0;
parameter W27TO35 = 0;
parameter W27TO36 = 0;
parameter W27TO37 = 0;
parameter W27TO38 = 0;
parameter W27TO39 = 0;
parameter W27TO40 = 0;
parameter W27TO41 = 0;
parameter W27TO42 = 0;
parameter W27TO43 = 0;
parameter W27TO44 = 0;
parameter W27TO45 = 0;
parameter W27TO46 = 0;
parameter W27TO47 = 0;
parameter W27TO48 = 0;
parameter W27TO49 = 0;
parameter W27TO50 = 0;
parameter W27TO51 = 0;
parameter W27TO52 = 0;
parameter W27TO53 = 0;
parameter W27TO54 = 0;
parameter W27TO55 = 0;
parameter W27TO56 = 0;
parameter W27TO57 = 0;
parameter W27TO58 = 0;
parameter W27TO59 = 0;
parameter W27TO60 = 0;
parameter W27TO61 = 0;
parameter W27TO62 = 0;
parameter W27TO63 = 0;
parameter W27TO64 = 0;
parameter W27TO65 = 0;
parameter W27TO66 = 0;
parameter W27TO67 = 0;
parameter W27TO68 = 0;
parameter W27TO69 = 0;
parameter W27TO70 = 0;
parameter W27TO71 = 0;
parameter W27TO72 = 0;
parameter W27TO73 = 0;
parameter W27TO74 = 0;
parameter W27TO75 = 0;
parameter W27TO76 = 0;
parameter W27TO77 = 0;
parameter W27TO78 = 0;
parameter W27TO79 = 0;
parameter W27TO80 = 0;
parameter W27TO81 = 0;
parameter W27TO82 = 0;
parameter W27TO83 = 0;
parameter W27TO84 = 0;
parameter W27TO85 = 0;
parameter W27TO86 = 0;
parameter W27TO87 = 0;
parameter W27TO88 = 0;
parameter W27TO89 = 0;
parameter W27TO90 = 0;
parameter W27TO91 = 0;
parameter W27TO92 = 0;
parameter W27TO93 = 0;
parameter W27TO94 = 0;
parameter W27TO95 = 0;
parameter W27TO96 = 0;
parameter W27TO97 = 0;
parameter W27TO98 = 0;
parameter W27TO99 = 0;
parameter W28TO0 = 0;
parameter W28TO1 = 0;
parameter W28TO2 = 0;
parameter W28TO3 = 0;
parameter W28TO4 = 0;
parameter W28TO5 = 0;
parameter W28TO6 = 0;
parameter W28TO7 = 0;
parameter W28TO8 = 0;
parameter W28TO9 = 0;
parameter W28TO10 = 0;
parameter W28TO11 = 0;
parameter W28TO12 = 0;
parameter W28TO13 = 0;
parameter W28TO14 = 0;
parameter W28TO15 = 0;
parameter W28TO16 = 0;
parameter W28TO17 = 0;
parameter W28TO18 = 0;
parameter W28TO19 = 0;
parameter W28TO20 = 0;
parameter W28TO21 = 0;
parameter W28TO22 = 0;
parameter W28TO23 = 0;
parameter W28TO24 = 0;
parameter W28TO25 = 0;
parameter W28TO26 = 0;
parameter W28TO27 = 0;
parameter W28TO28 = 0;
parameter W28TO29 = 0;
parameter W28TO30 = 0;
parameter W28TO31 = 0;
parameter W28TO32 = 0;
parameter W28TO33 = 0;
parameter W28TO34 = 0;
parameter W28TO35 = 0;
parameter W28TO36 = 0;
parameter W28TO37 = 0;
parameter W28TO38 = 0;
parameter W28TO39 = 0;
parameter W28TO40 = 0;
parameter W28TO41 = 0;
parameter W28TO42 = 0;
parameter W28TO43 = 0;
parameter W28TO44 = 0;
parameter W28TO45 = 0;
parameter W28TO46 = 0;
parameter W28TO47 = 0;
parameter W28TO48 = 0;
parameter W28TO49 = 0;
parameter W28TO50 = 0;
parameter W28TO51 = 0;
parameter W28TO52 = 0;
parameter W28TO53 = 0;
parameter W28TO54 = 0;
parameter W28TO55 = 0;
parameter W28TO56 = 0;
parameter W28TO57 = 0;
parameter W28TO58 = 0;
parameter W28TO59 = 0;
parameter W28TO60 = 0;
parameter W28TO61 = 0;
parameter W28TO62 = 0;
parameter W28TO63 = 0;
parameter W28TO64 = 0;
parameter W28TO65 = 0;
parameter W28TO66 = 0;
parameter W28TO67 = 0;
parameter W28TO68 = 0;
parameter W28TO69 = 0;
parameter W28TO70 = 0;
parameter W28TO71 = 0;
parameter W28TO72 = 0;
parameter W28TO73 = 0;
parameter W28TO74 = 0;
parameter W28TO75 = 0;
parameter W28TO76 = 0;
parameter W28TO77 = 0;
parameter W28TO78 = 0;
parameter W28TO79 = 0;
parameter W28TO80 = 0;
parameter W28TO81 = 0;
parameter W28TO82 = 0;
parameter W28TO83 = 0;
parameter W28TO84 = 0;
parameter W28TO85 = 0;
parameter W28TO86 = 0;
parameter W28TO87 = 0;
parameter W28TO88 = 0;
parameter W28TO89 = 0;
parameter W28TO90 = 0;
parameter W28TO91 = 0;
parameter W28TO92 = 0;
parameter W28TO93 = 0;
parameter W28TO94 = 0;
parameter W28TO95 = 0;
parameter W28TO96 = 0;
parameter W28TO97 = 0;
parameter W28TO98 = 0;
parameter W28TO99 = 0;
parameter W29TO0 = 0;
parameter W29TO1 = 0;
parameter W29TO2 = 0;
parameter W29TO3 = 0;
parameter W29TO4 = 0;
parameter W29TO5 = 0;
parameter W29TO6 = 0;
parameter W29TO7 = 0;
parameter W29TO8 = 0;
parameter W29TO9 = 0;
parameter W29TO10 = 0;
parameter W29TO11 = 0;
parameter W29TO12 = 0;
parameter W29TO13 = 0;
parameter W29TO14 = 0;
parameter W29TO15 = 0;
parameter W29TO16 = 0;
parameter W29TO17 = 0;
parameter W29TO18 = 0;
parameter W29TO19 = 0;
parameter W29TO20 = 0;
parameter W29TO21 = 0;
parameter W29TO22 = 0;
parameter W29TO23 = 0;
parameter W29TO24 = 0;
parameter W29TO25 = 0;
parameter W29TO26 = 0;
parameter W29TO27 = 0;
parameter W29TO28 = 0;
parameter W29TO29 = 0;
parameter W29TO30 = 0;
parameter W29TO31 = 0;
parameter W29TO32 = 0;
parameter W29TO33 = 0;
parameter W29TO34 = 0;
parameter W29TO35 = 0;
parameter W29TO36 = 0;
parameter W29TO37 = 0;
parameter W29TO38 = 0;
parameter W29TO39 = 0;
parameter W29TO40 = 0;
parameter W29TO41 = 0;
parameter W29TO42 = 0;
parameter W29TO43 = 0;
parameter W29TO44 = 0;
parameter W29TO45 = 0;
parameter W29TO46 = 0;
parameter W29TO47 = 0;
parameter W29TO48 = 0;
parameter W29TO49 = 0;
parameter W29TO50 = 0;
parameter W29TO51 = 0;
parameter W29TO52 = 0;
parameter W29TO53 = 0;
parameter W29TO54 = 0;
parameter W29TO55 = 0;
parameter W29TO56 = 0;
parameter W29TO57 = 0;
parameter W29TO58 = 0;
parameter W29TO59 = 0;
parameter W29TO60 = 0;
parameter W29TO61 = 0;
parameter W29TO62 = 0;
parameter W29TO63 = 0;
parameter W29TO64 = 0;
parameter W29TO65 = 0;
parameter W29TO66 = 0;
parameter W29TO67 = 0;
parameter W29TO68 = 0;
parameter W29TO69 = 0;
parameter W29TO70 = 0;
parameter W29TO71 = 0;
parameter W29TO72 = 0;
parameter W29TO73 = 0;
parameter W29TO74 = 0;
parameter W29TO75 = 0;
parameter W29TO76 = 0;
parameter W29TO77 = 0;
parameter W29TO78 = 0;
parameter W29TO79 = 0;
parameter W29TO80 = 0;
parameter W29TO81 = 0;
parameter W29TO82 = 0;
parameter W29TO83 = 0;
parameter W29TO84 = 0;
parameter W29TO85 = 0;
parameter W29TO86 = 0;
parameter W29TO87 = 0;
parameter W29TO88 = 0;
parameter W29TO89 = 0;
parameter W29TO90 = 0;
parameter W29TO91 = 0;
parameter W29TO92 = 0;
parameter W29TO93 = 0;
parameter W29TO94 = 0;
parameter W29TO95 = 0;
parameter W29TO96 = 0;
parameter W29TO97 = 0;
parameter W29TO98 = 0;
parameter W29TO99 = 0;
parameter W30TO0 = 0;
parameter W30TO1 = 0;
parameter W30TO2 = 0;
parameter W30TO3 = 0;
parameter W30TO4 = 0;
parameter W30TO5 = 0;
parameter W30TO6 = 0;
parameter W30TO7 = 0;
parameter W30TO8 = 0;
parameter W30TO9 = 0;
parameter W30TO10 = 0;
parameter W30TO11 = 0;
parameter W30TO12 = 0;
parameter W30TO13 = 0;
parameter W30TO14 = 0;
parameter W30TO15 = 0;
parameter W30TO16 = 0;
parameter W30TO17 = 0;
parameter W30TO18 = 0;
parameter W30TO19 = 0;
parameter W30TO20 = 0;
parameter W30TO21 = 0;
parameter W30TO22 = 0;
parameter W30TO23 = 0;
parameter W30TO24 = 0;
parameter W30TO25 = 0;
parameter W30TO26 = 0;
parameter W30TO27 = 0;
parameter W30TO28 = 0;
parameter W30TO29 = 0;
parameter W30TO30 = 0;
parameter W30TO31 = 0;
parameter W30TO32 = 0;
parameter W30TO33 = 0;
parameter W30TO34 = 0;
parameter W30TO35 = 0;
parameter W30TO36 = 0;
parameter W30TO37 = 0;
parameter W30TO38 = 0;
parameter W30TO39 = 0;
parameter W30TO40 = 0;
parameter W30TO41 = 0;
parameter W30TO42 = 0;
parameter W30TO43 = 0;
parameter W30TO44 = 0;
parameter W30TO45 = 0;
parameter W30TO46 = 0;
parameter W30TO47 = 0;
parameter W30TO48 = 0;
parameter W30TO49 = 0;
parameter W30TO50 = 0;
parameter W30TO51 = 0;
parameter W30TO52 = 0;
parameter W30TO53 = 0;
parameter W30TO54 = 0;
parameter W30TO55 = 0;
parameter W30TO56 = 0;
parameter W30TO57 = 0;
parameter W30TO58 = 0;
parameter W30TO59 = 0;
parameter W30TO60 = 0;
parameter W30TO61 = 0;
parameter W30TO62 = 0;
parameter W30TO63 = 0;
parameter W30TO64 = 0;
parameter W30TO65 = 0;
parameter W30TO66 = 0;
parameter W30TO67 = 0;
parameter W30TO68 = 0;
parameter W30TO69 = 0;
parameter W30TO70 = 0;
parameter W30TO71 = 0;
parameter W30TO72 = 0;
parameter W30TO73 = 0;
parameter W30TO74 = 0;
parameter W30TO75 = 0;
parameter W30TO76 = 0;
parameter W30TO77 = 0;
parameter W30TO78 = 0;
parameter W30TO79 = 0;
parameter W30TO80 = 0;
parameter W30TO81 = 0;
parameter W30TO82 = 0;
parameter W30TO83 = 0;
parameter W30TO84 = 0;
parameter W30TO85 = 0;
parameter W30TO86 = 0;
parameter W30TO87 = 0;
parameter W30TO88 = 0;
parameter W30TO89 = 0;
parameter W30TO90 = 0;
parameter W30TO91 = 0;
parameter W30TO92 = 0;
parameter W30TO93 = 0;
parameter W30TO94 = 0;
parameter W30TO95 = 0;
parameter W30TO96 = 0;
parameter W30TO97 = 0;
parameter W30TO98 = 0;
parameter W30TO99 = 0;
parameter W31TO0 = 0;
parameter W31TO1 = 0;
parameter W31TO2 = 0;
parameter W31TO3 = 0;
parameter W31TO4 = 0;
parameter W31TO5 = 0;
parameter W31TO6 = 0;
parameter W31TO7 = 0;
parameter W31TO8 = 0;
parameter W31TO9 = 0;
parameter W31TO10 = 0;
parameter W31TO11 = 0;
parameter W31TO12 = 0;
parameter W31TO13 = 0;
parameter W31TO14 = 0;
parameter W31TO15 = 0;
parameter W31TO16 = 0;
parameter W31TO17 = 0;
parameter W31TO18 = 0;
parameter W31TO19 = 0;
parameter W31TO20 = 0;
parameter W31TO21 = 0;
parameter W31TO22 = 0;
parameter W31TO23 = 0;
parameter W31TO24 = 0;
parameter W31TO25 = 0;
parameter W31TO26 = 0;
parameter W31TO27 = 0;
parameter W31TO28 = 0;
parameter W31TO29 = 0;
parameter W31TO30 = 0;
parameter W31TO31 = 0;
parameter W31TO32 = 0;
parameter W31TO33 = 0;
parameter W31TO34 = 0;
parameter W31TO35 = 0;
parameter W31TO36 = 0;
parameter W31TO37 = 0;
parameter W31TO38 = 0;
parameter W31TO39 = 0;
parameter W31TO40 = 0;
parameter W31TO41 = 0;
parameter W31TO42 = 0;
parameter W31TO43 = 0;
parameter W31TO44 = 0;
parameter W31TO45 = 0;
parameter W31TO46 = 0;
parameter W31TO47 = 0;
parameter W31TO48 = 0;
parameter W31TO49 = 0;
parameter W31TO50 = 0;
parameter W31TO51 = 0;
parameter W31TO52 = 0;
parameter W31TO53 = 0;
parameter W31TO54 = 0;
parameter W31TO55 = 0;
parameter W31TO56 = 0;
parameter W31TO57 = 0;
parameter W31TO58 = 0;
parameter W31TO59 = 0;
parameter W31TO60 = 0;
parameter W31TO61 = 0;
parameter W31TO62 = 0;
parameter W31TO63 = 0;
parameter W31TO64 = 0;
parameter W31TO65 = 0;
parameter W31TO66 = 0;
parameter W31TO67 = 0;
parameter W31TO68 = 0;
parameter W31TO69 = 0;
parameter W31TO70 = 0;
parameter W31TO71 = 0;
parameter W31TO72 = 0;
parameter W31TO73 = 0;
parameter W31TO74 = 0;
parameter W31TO75 = 0;
parameter W31TO76 = 0;
parameter W31TO77 = 0;
parameter W31TO78 = 0;
parameter W31TO79 = 0;
parameter W31TO80 = 0;
parameter W31TO81 = 0;
parameter W31TO82 = 0;
parameter W31TO83 = 0;
parameter W31TO84 = 0;
parameter W31TO85 = 0;
parameter W31TO86 = 0;
parameter W31TO87 = 0;
parameter W31TO88 = 0;
parameter W31TO89 = 0;
parameter W31TO90 = 0;
parameter W31TO91 = 0;
parameter W31TO92 = 0;
parameter W31TO93 = 0;
parameter W31TO94 = 0;
parameter W31TO95 = 0;
parameter W31TO96 = 0;
parameter W31TO97 = 0;
parameter W31TO98 = 0;
parameter W31TO99 = 0;
parameter W32TO0 = 0;
parameter W32TO1 = 0;
parameter W32TO2 = 0;
parameter W32TO3 = 0;
parameter W32TO4 = 0;
parameter W32TO5 = 0;
parameter W32TO6 = 0;
parameter W32TO7 = 0;
parameter W32TO8 = 0;
parameter W32TO9 = 0;
parameter W32TO10 = 0;
parameter W32TO11 = 0;
parameter W32TO12 = 0;
parameter W32TO13 = 0;
parameter W32TO14 = 0;
parameter W32TO15 = 0;
parameter W32TO16 = 0;
parameter W32TO17 = 0;
parameter W32TO18 = 0;
parameter W32TO19 = 0;
parameter W32TO20 = 0;
parameter W32TO21 = 0;
parameter W32TO22 = 0;
parameter W32TO23 = 0;
parameter W32TO24 = 0;
parameter W32TO25 = 0;
parameter W32TO26 = 0;
parameter W32TO27 = 0;
parameter W32TO28 = 0;
parameter W32TO29 = 0;
parameter W32TO30 = 0;
parameter W32TO31 = 0;
parameter W32TO32 = 0;
parameter W32TO33 = 0;
parameter W32TO34 = 0;
parameter W32TO35 = 0;
parameter W32TO36 = 0;
parameter W32TO37 = 0;
parameter W32TO38 = 0;
parameter W32TO39 = 0;
parameter W32TO40 = 0;
parameter W32TO41 = 0;
parameter W32TO42 = 0;
parameter W32TO43 = 0;
parameter W32TO44 = 0;
parameter W32TO45 = 0;
parameter W32TO46 = 0;
parameter W32TO47 = 0;
parameter W32TO48 = 0;
parameter W32TO49 = 0;
parameter W32TO50 = 0;
parameter W32TO51 = 0;
parameter W32TO52 = 0;
parameter W32TO53 = 0;
parameter W32TO54 = 0;
parameter W32TO55 = 0;
parameter W32TO56 = 0;
parameter W32TO57 = 0;
parameter W32TO58 = 0;
parameter W32TO59 = 0;
parameter W32TO60 = 0;
parameter W32TO61 = 0;
parameter W32TO62 = 0;
parameter W32TO63 = 0;
parameter W32TO64 = 0;
parameter W32TO65 = 0;
parameter W32TO66 = 0;
parameter W32TO67 = 0;
parameter W32TO68 = 0;
parameter W32TO69 = 0;
parameter W32TO70 = 0;
parameter W32TO71 = 0;
parameter W32TO72 = 0;
parameter W32TO73 = 0;
parameter W32TO74 = 0;
parameter W32TO75 = 0;
parameter W32TO76 = 0;
parameter W32TO77 = 0;
parameter W32TO78 = 0;
parameter W32TO79 = 0;
parameter W32TO80 = 0;
parameter W32TO81 = 0;
parameter W32TO82 = 0;
parameter W32TO83 = 0;
parameter W32TO84 = 0;
parameter W32TO85 = 0;
parameter W32TO86 = 0;
parameter W32TO87 = 0;
parameter W32TO88 = 0;
parameter W32TO89 = 0;
parameter W32TO90 = 0;
parameter W32TO91 = 0;
parameter W32TO92 = 0;
parameter W32TO93 = 0;
parameter W32TO94 = 0;
parameter W32TO95 = 0;
parameter W32TO96 = 0;
parameter W32TO97 = 0;
parameter W32TO98 = 0;
parameter W32TO99 = 0;
parameter W33TO0 = 0;
parameter W33TO1 = 0;
parameter W33TO2 = 0;
parameter W33TO3 = 0;
parameter W33TO4 = 0;
parameter W33TO5 = 0;
parameter W33TO6 = 0;
parameter W33TO7 = 0;
parameter W33TO8 = 0;
parameter W33TO9 = 0;
parameter W33TO10 = 0;
parameter W33TO11 = 0;
parameter W33TO12 = 0;
parameter W33TO13 = 0;
parameter W33TO14 = 0;
parameter W33TO15 = 0;
parameter W33TO16 = 0;
parameter W33TO17 = 0;
parameter W33TO18 = 0;
parameter W33TO19 = 0;
parameter W33TO20 = 0;
parameter W33TO21 = 0;
parameter W33TO22 = 0;
parameter W33TO23 = 0;
parameter W33TO24 = 0;
parameter W33TO25 = 0;
parameter W33TO26 = 0;
parameter W33TO27 = 0;
parameter W33TO28 = 0;
parameter W33TO29 = 0;
parameter W33TO30 = 0;
parameter W33TO31 = 0;
parameter W33TO32 = 0;
parameter W33TO33 = 0;
parameter W33TO34 = 0;
parameter W33TO35 = 0;
parameter W33TO36 = 0;
parameter W33TO37 = 0;
parameter W33TO38 = 0;
parameter W33TO39 = 0;
parameter W33TO40 = 0;
parameter W33TO41 = 0;
parameter W33TO42 = 0;
parameter W33TO43 = 0;
parameter W33TO44 = 0;
parameter W33TO45 = 0;
parameter W33TO46 = 0;
parameter W33TO47 = 0;
parameter W33TO48 = 0;
parameter W33TO49 = 0;
parameter W33TO50 = 0;
parameter W33TO51 = 0;
parameter W33TO52 = 0;
parameter W33TO53 = 0;
parameter W33TO54 = 0;
parameter W33TO55 = 0;
parameter W33TO56 = 0;
parameter W33TO57 = 0;
parameter W33TO58 = 0;
parameter W33TO59 = 0;
parameter W33TO60 = 0;
parameter W33TO61 = 0;
parameter W33TO62 = 0;
parameter W33TO63 = 0;
parameter W33TO64 = 0;
parameter W33TO65 = 0;
parameter W33TO66 = 0;
parameter W33TO67 = 0;
parameter W33TO68 = 0;
parameter W33TO69 = 0;
parameter W33TO70 = 0;
parameter W33TO71 = 0;
parameter W33TO72 = 0;
parameter W33TO73 = 0;
parameter W33TO74 = 0;
parameter W33TO75 = 0;
parameter W33TO76 = 0;
parameter W33TO77 = 0;
parameter W33TO78 = 0;
parameter W33TO79 = 0;
parameter W33TO80 = 0;
parameter W33TO81 = 0;
parameter W33TO82 = 0;
parameter W33TO83 = 0;
parameter W33TO84 = 0;
parameter W33TO85 = 0;
parameter W33TO86 = 0;
parameter W33TO87 = 0;
parameter W33TO88 = 0;
parameter W33TO89 = 0;
parameter W33TO90 = 0;
parameter W33TO91 = 0;
parameter W33TO92 = 0;
parameter W33TO93 = 0;
parameter W33TO94 = 0;
parameter W33TO95 = 0;
parameter W33TO96 = 0;
parameter W33TO97 = 0;
parameter W33TO98 = 0;
parameter W33TO99 = 0;
parameter W34TO0 = 0;
parameter W34TO1 = 0;
parameter W34TO2 = 0;
parameter W34TO3 = 0;
parameter W34TO4 = 0;
parameter W34TO5 = 0;
parameter W34TO6 = 0;
parameter W34TO7 = 0;
parameter W34TO8 = 0;
parameter W34TO9 = 0;
parameter W34TO10 = 0;
parameter W34TO11 = 0;
parameter W34TO12 = 0;
parameter W34TO13 = 0;
parameter W34TO14 = 0;
parameter W34TO15 = 0;
parameter W34TO16 = 0;
parameter W34TO17 = 0;
parameter W34TO18 = 0;
parameter W34TO19 = 0;
parameter W34TO20 = 0;
parameter W34TO21 = 0;
parameter W34TO22 = 0;
parameter W34TO23 = 0;
parameter W34TO24 = 0;
parameter W34TO25 = 0;
parameter W34TO26 = 0;
parameter W34TO27 = 0;
parameter W34TO28 = 0;
parameter W34TO29 = 0;
parameter W34TO30 = 0;
parameter W34TO31 = 0;
parameter W34TO32 = 0;
parameter W34TO33 = 0;
parameter W34TO34 = 0;
parameter W34TO35 = 0;
parameter W34TO36 = 0;
parameter W34TO37 = 0;
parameter W34TO38 = 0;
parameter W34TO39 = 0;
parameter W34TO40 = 0;
parameter W34TO41 = 0;
parameter W34TO42 = 0;
parameter W34TO43 = 0;
parameter W34TO44 = 0;
parameter W34TO45 = 0;
parameter W34TO46 = 0;
parameter W34TO47 = 0;
parameter W34TO48 = 0;
parameter W34TO49 = 0;
parameter W34TO50 = 0;
parameter W34TO51 = 0;
parameter W34TO52 = 0;
parameter W34TO53 = 0;
parameter W34TO54 = 0;
parameter W34TO55 = 0;
parameter W34TO56 = 0;
parameter W34TO57 = 0;
parameter W34TO58 = 0;
parameter W34TO59 = 0;
parameter W34TO60 = 0;
parameter W34TO61 = 0;
parameter W34TO62 = 0;
parameter W34TO63 = 0;
parameter W34TO64 = 0;
parameter W34TO65 = 0;
parameter W34TO66 = 0;
parameter W34TO67 = 0;
parameter W34TO68 = 0;
parameter W34TO69 = 0;
parameter W34TO70 = 0;
parameter W34TO71 = 0;
parameter W34TO72 = 0;
parameter W34TO73 = 0;
parameter W34TO74 = 0;
parameter W34TO75 = 0;
parameter W34TO76 = 0;
parameter W34TO77 = 0;
parameter W34TO78 = 0;
parameter W34TO79 = 0;
parameter W34TO80 = 0;
parameter W34TO81 = 0;
parameter W34TO82 = 0;
parameter W34TO83 = 0;
parameter W34TO84 = 0;
parameter W34TO85 = 0;
parameter W34TO86 = 0;
parameter W34TO87 = 0;
parameter W34TO88 = 0;
parameter W34TO89 = 0;
parameter W34TO90 = 0;
parameter W34TO91 = 0;
parameter W34TO92 = 0;
parameter W34TO93 = 0;
parameter W34TO94 = 0;
parameter W34TO95 = 0;
parameter W34TO96 = 0;
parameter W34TO97 = 0;
parameter W34TO98 = 0;
parameter W34TO99 = 0;
parameter W35TO0 = 0;
parameter W35TO1 = 0;
parameter W35TO2 = 0;
parameter W35TO3 = 0;
parameter W35TO4 = 0;
parameter W35TO5 = 0;
parameter W35TO6 = 0;
parameter W35TO7 = 0;
parameter W35TO8 = 0;
parameter W35TO9 = 0;
parameter W35TO10 = 0;
parameter W35TO11 = 0;
parameter W35TO12 = 0;
parameter W35TO13 = 0;
parameter W35TO14 = 0;
parameter W35TO15 = 0;
parameter W35TO16 = 0;
parameter W35TO17 = 0;
parameter W35TO18 = 0;
parameter W35TO19 = 0;
parameter W35TO20 = 0;
parameter W35TO21 = 0;
parameter W35TO22 = 0;
parameter W35TO23 = 0;
parameter W35TO24 = 0;
parameter W35TO25 = 0;
parameter W35TO26 = 0;
parameter W35TO27 = 0;
parameter W35TO28 = 0;
parameter W35TO29 = 0;
parameter W35TO30 = 0;
parameter W35TO31 = 0;
parameter W35TO32 = 0;
parameter W35TO33 = 0;
parameter W35TO34 = 0;
parameter W35TO35 = 0;
parameter W35TO36 = 0;
parameter W35TO37 = 0;
parameter W35TO38 = 0;
parameter W35TO39 = 0;
parameter W35TO40 = 0;
parameter W35TO41 = 0;
parameter W35TO42 = 0;
parameter W35TO43 = 0;
parameter W35TO44 = 0;
parameter W35TO45 = 0;
parameter W35TO46 = 0;
parameter W35TO47 = 0;
parameter W35TO48 = 0;
parameter W35TO49 = 0;
parameter W35TO50 = 0;
parameter W35TO51 = 0;
parameter W35TO52 = 0;
parameter W35TO53 = 0;
parameter W35TO54 = 0;
parameter W35TO55 = 0;
parameter W35TO56 = 0;
parameter W35TO57 = 0;
parameter W35TO58 = 0;
parameter W35TO59 = 0;
parameter W35TO60 = 0;
parameter W35TO61 = 0;
parameter W35TO62 = 0;
parameter W35TO63 = 0;
parameter W35TO64 = 0;
parameter W35TO65 = 0;
parameter W35TO66 = 0;
parameter W35TO67 = 0;
parameter W35TO68 = 0;
parameter W35TO69 = 0;
parameter W35TO70 = 0;
parameter W35TO71 = 0;
parameter W35TO72 = 0;
parameter W35TO73 = 0;
parameter W35TO74 = 0;
parameter W35TO75 = 0;
parameter W35TO76 = 0;
parameter W35TO77 = 0;
parameter W35TO78 = 0;
parameter W35TO79 = 0;
parameter W35TO80 = 0;
parameter W35TO81 = 0;
parameter W35TO82 = 0;
parameter W35TO83 = 0;
parameter W35TO84 = 0;
parameter W35TO85 = 0;
parameter W35TO86 = 0;
parameter W35TO87 = 0;
parameter W35TO88 = 0;
parameter W35TO89 = 0;
parameter W35TO90 = 0;
parameter W35TO91 = 0;
parameter W35TO92 = 0;
parameter W35TO93 = 0;
parameter W35TO94 = 0;
parameter W35TO95 = 0;
parameter W35TO96 = 0;
parameter W35TO97 = 0;
parameter W35TO98 = 0;
parameter W35TO99 = 0;
parameter W36TO0 = 0;
parameter W36TO1 = 0;
parameter W36TO2 = 0;
parameter W36TO3 = 0;
parameter W36TO4 = 0;
parameter W36TO5 = 0;
parameter W36TO6 = 0;
parameter W36TO7 = 0;
parameter W36TO8 = 0;
parameter W36TO9 = 0;
parameter W36TO10 = 0;
parameter W36TO11 = 0;
parameter W36TO12 = 0;
parameter W36TO13 = 0;
parameter W36TO14 = 0;
parameter W36TO15 = 0;
parameter W36TO16 = 0;
parameter W36TO17 = 0;
parameter W36TO18 = 0;
parameter W36TO19 = 0;
parameter W36TO20 = 0;
parameter W36TO21 = 0;
parameter W36TO22 = 0;
parameter W36TO23 = 0;
parameter W36TO24 = 0;
parameter W36TO25 = 0;
parameter W36TO26 = 0;
parameter W36TO27 = 0;
parameter W36TO28 = 0;
parameter W36TO29 = 0;
parameter W36TO30 = 0;
parameter W36TO31 = 0;
parameter W36TO32 = 0;
parameter W36TO33 = 0;
parameter W36TO34 = 0;
parameter W36TO35 = 0;
parameter W36TO36 = 0;
parameter W36TO37 = 0;
parameter W36TO38 = 0;
parameter W36TO39 = 0;
parameter W36TO40 = 0;
parameter W36TO41 = 0;
parameter W36TO42 = 0;
parameter W36TO43 = 0;
parameter W36TO44 = 0;
parameter W36TO45 = 0;
parameter W36TO46 = 0;
parameter W36TO47 = 0;
parameter W36TO48 = 0;
parameter W36TO49 = 0;
parameter W36TO50 = 0;
parameter W36TO51 = 0;
parameter W36TO52 = 0;
parameter W36TO53 = 0;
parameter W36TO54 = 0;
parameter W36TO55 = 0;
parameter W36TO56 = 0;
parameter W36TO57 = 0;
parameter W36TO58 = 0;
parameter W36TO59 = 0;
parameter W36TO60 = 0;
parameter W36TO61 = 0;
parameter W36TO62 = 0;
parameter W36TO63 = 0;
parameter W36TO64 = 0;
parameter W36TO65 = 0;
parameter W36TO66 = 0;
parameter W36TO67 = 0;
parameter W36TO68 = 0;
parameter W36TO69 = 0;
parameter W36TO70 = 0;
parameter W36TO71 = 0;
parameter W36TO72 = 0;
parameter W36TO73 = 0;
parameter W36TO74 = 0;
parameter W36TO75 = 0;
parameter W36TO76 = 0;
parameter W36TO77 = 0;
parameter W36TO78 = 0;
parameter W36TO79 = 0;
parameter W36TO80 = 0;
parameter W36TO81 = 0;
parameter W36TO82 = 0;
parameter W36TO83 = 0;
parameter W36TO84 = 0;
parameter W36TO85 = 0;
parameter W36TO86 = 0;
parameter W36TO87 = 0;
parameter W36TO88 = 0;
parameter W36TO89 = 0;
parameter W36TO90 = 0;
parameter W36TO91 = 0;
parameter W36TO92 = 0;
parameter W36TO93 = 0;
parameter W36TO94 = 0;
parameter W36TO95 = 0;
parameter W36TO96 = 0;
parameter W36TO97 = 0;
parameter W36TO98 = 0;
parameter W36TO99 = 0;
parameter W37TO0 = 0;
parameter W37TO1 = 0;
parameter W37TO2 = 0;
parameter W37TO3 = 0;
parameter W37TO4 = 0;
parameter W37TO5 = 0;
parameter W37TO6 = 0;
parameter W37TO7 = 0;
parameter W37TO8 = 0;
parameter W37TO9 = 0;
parameter W37TO10 = 0;
parameter W37TO11 = 0;
parameter W37TO12 = 0;
parameter W37TO13 = 0;
parameter W37TO14 = 0;
parameter W37TO15 = 0;
parameter W37TO16 = 0;
parameter W37TO17 = 0;
parameter W37TO18 = 0;
parameter W37TO19 = 0;
parameter W37TO20 = 0;
parameter W37TO21 = 0;
parameter W37TO22 = 0;
parameter W37TO23 = 0;
parameter W37TO24 = 0;
parameter W37TO25 = 0;
parameter W37TO26 = 0;
parameter W37TO27 = 0;
parameter W37TO28 = 0;
parameter W37TO29 = 0;
parameter W37TO30 = 0;
parameter W37TO31 = 0;
parameter W37TO32 = 0;
parameter W37TO33 = 0;
parameter W37TO34 = 0;
parameter W37TO35 = 0;
parameter W37TO36 = 0;
parameter W37TO37 = 0;
parameter W37TO38 = 0;
parameter W37TO39 = 0;
parameter W37TO40 = 0;
parameter W37TO41 = 0;
parameter W37TO42 = 0;
parameter W37TO43 = 0;
parameter W37TO44 = 0;
parameter W37TO45 = 0;
parameter W37TO46 = 0;
parameter W37TO47 = 0;
parameter W37TO48 = 0;
parameter W37TO49 = 0;
parameter W37TO50 = 0;
parameter W37TO51 = 0;
parameter W37TO52 = 0;
parameter W37TO53 = 0;
parameter W37TO54 = 0;
parameter W37TO55 = 0;
parameter W37TO56 = 0;
parameter W37TO57 = 0;
parameter W37TO58 = 0;
parameter W37TO59 = 0;
parameter W37TO60 = 0;
parameter W37TO61 = 0;
parameter W37TO62 = 0;
parameter W37TO63 = 0;
parameter W37TO64 = 0;
parameter W37TO65 = 0;
parameter W37TO66 = 0;
parameter W37TO67 = 0;
parameter W37TO68 = 0;
parameter W37TO69 = 0;
parameter W37TO70 = 0;
parameter W37TO71 = 0;
parameter W37TO72 = 0;
parameter W37TO73 = 0;
parameter W37TO74 = 0;
parameter W37TO75 = 0;
parameter W37TO76 = 0;
parameter W37TO77 = 0;
parameter W37TO78 = 0;
parameter W37TO79 = 0;
parameter W37TO80 = 0;
parameter W37TO81 = 0;
parameter W37TO82 = 0;
parameter W37TO83 = 0;
parameter W37TO84 = 0;
parameter W37TO85 = 0;
parameter W37TO86 = 0;
parameter W37TO87 = 0;
parameter W37TO88 = 0;
parameter W37TO89 = 0;
parameter W37TO90 = 0;
parameter W37TO91 = 0;
parameter W37TO92 = 0;
parameter W37TO93 = 0;
parameter W37TO94 = 0;
parameter W37TO95 = 0;
parameter W37TO96 = 0;
parameter W37TO97 = 0;
parameter W37TO98 = 0;
parameter W37TO99 = 0;
parameter W38TO0 = 0;
parameter W38TO1 = 0;
parameter W38TO2 = 0;
parameter W38TO3 = 0;
parameter W38TO4 = 0;
parameter W38TO5 = 0;
parameter W38TO6 = 0;
parameter W38TO7 = 0;
parameter W38TO8 = 0;
parameter W38TO9 = 0;
parameter W38TO10 = 0;
parameter W38TO11 = 0;
parameter W38TO12 = 0;
parameter W38TO13 = 0;
parameter W38TO14 = 0;
parameter W38TO15 = 0;
parameter W38TO16 = 0;
parameter W38TO17 = 0;
parameter W38TO18 = 0;
parameter W38TO19 = 0;
parameter W38TO20 = 0;
parameter W38TO21 = 0;
parameter W38TO22 = 0;
parameter W38TO23 = 0;
parameter W38TO24 = 0;
parameter W38TO25 = 0;
parameter W38TO26 = 0;
parameter W38TO27 = 0;
parameter W38TO28 = 0;
parameter W38TO29 = 0;
parameter W38TO30 = 0;
parameter W38TO31 = 0;
parameter W38TO32 = 0;
parameter W38TO33 = 0;
parameter W38TO34 = 0;
parameter W38TO35 = 0;
parameter W38TO36 = 0;
parameter W38TO37 = 0;
parameter W38TO38 = 0;
parameter W38TO39 = 0;
parameter W38TO40 = 0;
parameter W38TO41 = 0;
parameter W38TO42 = 0;
parameter W38TO43 = 0;
parameter W38TO44 = 0;
parameter W38TO45 = 0;
parameter W38TO46 = 0;
parameter W38TO47 = 0;
parameter W38TO48 = 0;
parameter W38TO49 = 0;
parameter W38TO50 = 0;
parameter W38TO51 = 0;
parameter W38TO52 = 0;
parameter W38TO53 = 0;
parameter W38TO54 = 0;
parameter W38TO55 = 0;
parameter W38TO56 = 0;
parameter W38TO57 = 0;
parameter W38TO58 = 0;
parameter W38TO59 = 0;
parameter W38TO60 = 0;
parameter W38TO61 = 0;
parameter W38TO62 = 0;
parameter W38TO63 = 0;
parameter W38TO64 = 0;
parameter W38TO65 = 0;
parameter W38TO66 = 0;
parameter W38TO67 = 0;
parameter W38TO68 = 0;
parameter W38TO69 = 0;
parameter W38TO70 = 0;
parameter W38TO71 = 0;
parameter W38TO72 = 0;
parameter W38TO73 = 0;
parameter W38TO74 = 0;
parameter W38TO75 = 0;
parameter W38TO76 = 0;
parameter W38TO77 = 0;
parameter W38TO78 = 0;
parameter W38TO79 = 0;
parameter W38TO80 = 0;
parameter W38TO81 = 0;
parameter W38TO82 = 0;
parameter W38TO83 = 0;
parameter W38TO84 = 0;
parameter W38TO85 = 0;
parameter W38TO86 = 0;
parameter W38TO87 = 0;
parameter W38TO88 = 0;
parameter W38TO89 = 0;
parameter W38TO90 = 0;
parameter W38TO91 = 0;
parameter W38TO92 = 0;
parameter W38TO93 = 0;
parameter W38TO94 = 0;
parameter W38TO95 = 0;
parameter W38TO96 = 0;
parameter W38TO97 = 0;
parameter W38TO98 = 0;
parameter W38TO99 = 0;
parameter W39TO0 = 0;
parameter W39TO1 = 0;
parameter W39TO2 = 0;
parameter W39TO3 = 0;
parameter W39TO4 = 0;
parameter W39TO5 = 0;
parameter W39TO6 = 0;
parameter W39TO7 = 0;
parameter W39TO8 = 0;
parameter W39TO9 = 0;
parameter W39TO10 = 0;
parameter W39TO11 = 0;
parameter W39TO12 = 0;
parameter W39TO13 = 0;
parameter W39TO14 = 0;
parameter W39TO15 = 0;
parameter W39TO16 = 0;
parameter W39TO17 = 0;
parameter W39TO18 = 0;
parameter W39TO19 = 0;
parameter W39TO20 = 0;
parameter W39TO21 = 0;
parameter W39TO22 = 0;
parameter W39TO23 = 0;
parameter W39TO24 = 0;
parameter W39TO25 = 0;
parameter W39TO26 = 0;
parameter W39TO27 = 0;
parameter W39TO28 = 0;
parameter W39TO29 = 0;
parameter W39TO30 = 0;
parameter W39TO31 = 0;
parameter W39TO32 = 0;
parameter W39TO33 = 0;
parameter W39TO34 = 0;
parameter W39TO35 = 0;
parameter W39TO36 = 0;
parameter W39TO37 = 0;
parameter W39TO38 = 0;
parameter W39TO39 = 0;
parameter W39TO40 = 0;
parameter W39TO41 = 0;
parameter W39TO42 = 0;
parameter W39TO43 = 0;
parameter W39TO44 = 0;
parameter W39TO45 = 0;
parameter W39TO46 = 0;
parameter W39TO47 = 0;
parameter W39TO48 = 0;
parameter W39TO49 = 0;
parameter W39TO50 = 0;
parameter W39TO51 = 0;
parameter W39TO52 = 0;
parameter W39TO53 = 0;
parameter W39TO54 = 0;
parameter W39TO55 = 0;
parameter W39TO56 = 0;
parameter W39TO57 = 0;
parameter W39TO58 = 0;
parameter W39TO59 = 0;
parameter W39TO60 = 0;
parameter W39TO61 = 0;
parameter W39TO62 = 0;
parameter W39TO63 = 0;
parameter W39TO64 = 0;
parameter W39TO65 = 0;
parameter W39TO66 = 0;
parameter W39TO67 = 0;
parameter W39TO68 = 0;
parameter W39TO69 = 0;
parameter W39TO70 = 0;
parameter W39TO71 = 0;
parameter W39TO72 = 0;
parameter W39TO73 = 0;
parameter W39TO74 = 0;
parameter W39TO75 = 0;
parameter W39TO76 = 0;
parameter W39TO77 = 0;
parameter W39TO78 = 0;
parameter W39TO79 = 0;
parameter W39TO80 = 0;
parameter W39TO81 = 0;
parameter W39TO82 = 0;
parameter W39TO83 = 0;
parameter W39TO84 = 0;
parameter W39TO85 = 0;
parameter W39TO86 = 0;
parameter W39TO87 = 0;
parameter W39TO88 = 0;
parameter W39TO89 = 0;
parameter W39TO90 = 0;
parameter W39TO91 = 0;
parameter W39TO92 = 0;
parameter W39TO93 = 0;
parameter W39TO94 = 0;
parameter W39TO95 = 0;
parameter W39TO96 = 0;
parameter W39TO97 = 0;
parameter W39TO98 = 0;
parameter W39TO99 = 0;
parameter W40TO0 = 0;
parameter W40TO1 = 0;
parameter W40TO2 = 0;
parameter W40TO3 = 0;
parameter W40TO4 = 0;
parameter W40TO5 = 0;
parameter W40TO6 = 0;
parameter W40TO7 = 0;
parameter W40TO8 = 0;
parameter W40TO9 = 0;
parameter W40TO10 = 0;
parameter W40TO11 = 0;
parameter W40TO12 = 0;
parameter W40TO13 = 0;
parameter W40TO14 = 0;
parameter W40TO15 = 0;
parameter W40TO16 = 0;
parameter W40TO17 = 0;
parameter W40TO18 = 0;
parameter W40TO19 = 0;
parameter W40TO20 = 0;
parameter W40TO21 = 0;
parameter W40TO22 = 0;
parameter W40TO23 = 0;
parameter W40TO24 = 0;
parameter W40TO25 = 0;
parameter W40TO26 = 0;
parameter W40TO27 = 0;
parameter W40TO28 = 0;
parameter W40TO29 = 0;
parameter W40TO30 = 0;
parameter W40TO31 = 0;
parameter W40TO32 = 0;
parameter W40TO33 = 0;
parameter W40TO34 = 0;
parameter W40TO35 = 0;
parameter W40TO36 = 0;
parameter W40TO37 = 0;
parameter W40TO38 = 0;
parameter W40TO39 = 0;
parameter W40TO40 = 0;
parameter W40TO41 = 0;
parameter W40TO42 = 0;
parameter W40TO43 = 0;
parameter W40TO44 = 0;
parameter W40TO45 = 0;
parameter W40TO46 = 0;
parameter W40TO47 = 0;
parameter W40TO48 = 0;
parameter W40TO49 = 0;
parameter W40TO50 = 0;
parameter W40TO51 = 0;
parameter W40TO52 = 0;
parameter W40TO53 = 0;
parameter W40TO54 = 0;
parameter W40TO55 = 0;
parameter W40TO56 = 0;
parameter W40TO57 = 0;
parameter W40TO58 = 0;
parameter W40TO59 = 0;
parameter W40TO60 = 0;
parameter W40TO61 = 0;
parameter W40TO62 = 0;
parameter W40TO63 = 0;
parameter W40TO64 = 0;
parameter W40TO65 = 0;
parameter W40TO66 = 0;
parameter W40TO67 = 0;
parameter W40TO68 = 0;
parameter W40TO69 = 0;
parameter W40TO70 = 0;
parameter W40TO71 = 0;
parameter W40TO72 = 0;
parameter W40TO73 = 0;
parameter W40TO74 = 0;
parameter W40TO75 = 0;
parameter W40TO76 = 0;
parameter W40TO77 = 0;
parameter W40TO78 = 0;
parameter W40TO79 = 0;
parameter W40TO80 = 0;
parameter W40TO81 = 0;
parameter W40TO82 = 0;
parameter W40TO83 = 0;
parameter W40TO84 = 0;
parameter W40TO85 = 0;
parameter W40TO86 = 0;
parameter W40TO87 = 0;
parameter W40TO88 = 0;
parameter W40TO89 = 0;
parameter W40TO90 = 0;
parameter W40TO91 = 0;
parameter W40TO92 = 0;
parameter W40TO93 = 0;
parameter W40TO94 = 0;
parameter W40TO95 = 0;
parameter W40TO96 = 0;
parameter W40TO97 = 0;
parameter W40TO98 = 0;
parameter W40TO99 = 0;
parameter W41TO0 = 0;
parameter W41TO1 = 0;
parameter W41TO2 = 0;
parameter W41TO3 = 0;
parameter W41TO4 = 0;
parameter W41TO5 = 0;
parameter W41TO6 = 0;
parameter W41TO7 = 0;
parameter W41TO8 = 0;
parameter W41TO9 = 0;
parameter W41TO10 = 0;
parameter W41TO11 = 0;
parameter W41TO12 = 0;
parameter W41TO13 = 0;
parameter W41TO14 = 0;
parameter W41TO15 = 0;
parameter W41TO16 = 0;
parameter W41TO17 = 0;
parameter W41TO18 = 0;
parameter W41TO19 = 0;
parameter W41TO20 = 0;
parameter W41TO21 = 0;
parameter W41TO22 = 0;
parameter W41TO23 = 0;
parameter W41TO24 = 0;
parameter W41TO25 = 0;
parameter W41TO26 = 0;
parameter W41TO27 = 0;
parameter W41TO28 = 0;
parameter W41TO29 = 0;
parameter W41TO30 = 0;
parameter W41TO31 = 0;
parameter W41TO32 = 0;
parameter W41TO33 = 0;
parameter W41TO34 = 0;
parameter W41TO35 = 0;
parameter W41TO36 = 0;
parameter W41TO37 = 0;
parameter W41TO38 = 0;
parameter W41TO39 = 0;
parameter W41TO40 = 0;
parameter W41TO41 = 0;
parameter W41TO42 = 0;
parameter W41TO43 = 0;
parameter W41TO44 = 0;
parameter W41TO45 = 0;
parameter W41TO46 = 0;
parameter W41TO47 = 0;
parameter W41TO48 = 0;
parameter W41TO49 = 0;
parameter W41TO50 = 0;
parameter W41TO51 = 0;
parameter W41TO52 = 0;
parameter W41TO53 = 0;
parameter W41TO54 = 0;
parameter W41TO55 = 0;
parameter W41TO56 = 0;
parameter W41TO57 = 0;
parameter W41TO58 = 0;
parameter W41TO59 = 0;
parameter W41TO60 = 0;
parameter W41TO61 = 0;
parameter W41TO62 = 0;
parameter W41TO63 = 0;
parameter W41TO64 = 0;
parameter W41TO65 = 0;
parameter W41TO66 = 0;
parameter W41TO67 = 0;
parameter W41TO68 = 0;
parameter W41TO69 = 0;
parameter W41TO70 = 0;
parameter W41TO71 = 0;
parameter W41TO72 = 0;
parameter W41TO73 = 0;
parameter W41TO74 = 0;
parameter W41TO75 = 0;
parameter W41TO76 = 0;
parameter W41TO77 = 0;
parameter W41TO78 = 0;
parameter W41TO79 = 0;
parameter W41TO80 = 0;
parameter W41TO81 = 0;
parameter W41TO82 = 0;
parameter W41TO83 = 0;
parameter W41TO84 = 0;
parameter W41TO85 = 0;
parameter W41TO86 = 0;
parameter W41TO87 = 0;
parameter W41TO88 = 0;
parameter W41TO89 = 0;
parameter W41TO90 = 0;
parameter W41TO91 = 0;
parameter W41TO92 = 0;
parameter W41TO93 = 0;
parameter W41TO94 = 0;
parameter W41TO95 = 0;
parameter W41TO96 = 0;
parameter W41TO97 = 0;
parameter W41TO98 = 0;
parameter W41TO99 = 0;
parameter W42TO0 = 0;
parameter W42TO1 = 0;
parameter W42TO2 = 0;
parameter W42TO3 = 0;
parameter W42TO4 = 0;
parameter W42TO5 = 0;
parameter W42TO6 = 0;
parameter W42TO7 = 0;
parameter W42TO8 = 0;
parameter W42TO9 = 0;
parameter W42TO10 = 0;
parameter W42TO11 = 0;
parameter W42TO12 = 0;
parameter W42TO13 = 0;
parameter W42TO14 = 0;
parameter W42TO15 = 0;
parameter W42TO16 = 0;
parameter W42TO17 = 0;
parameter W42TO18 = 0;
parameter W42TO19 = 0;
parameter W42TO20 = 0;
parameter W42TO21 = 0;
parameter W42TO22 = 0;
parameter W42TO23 = 0;
parameter W42TO24 = 0;
parameter W42TO25 = 0;
parameter W42TO26 = 0;
parameter W42TO27 = 0;
parameter W42TO28 = 0;
parameter W42TO29 = 0;
parameter W42TO30 = 0;
parameter W42TO31 = 0;
parameter W42TO32 = 0;
parameter W42TO33 = 0;
parameter W42TO34 = 0;
parameter W42TO35 = 0;
parameter W42TO36 = 0;
parameter W42TO37 = 0;
parameter W42TO38 = 0;
parameter W42TO39 = 0;
parameter W42TO40 = 0;
parameter W42TO41 = 0;
parameter W42TO42 = 0;
parameter W42TO43 = 0;
parameter W42TO44 = 0;
parameter W42TO45 = 0;
parameter W42TO46 = 0;
parameter W42TO47 = 0;
parameter W42TO48 = 0;
parameter W42TO49 = 0;
parameter W42TO50 = 0;
parameter W42TO51 = 0;
parameter W42TO52 = 0;
parameter W42TO53 = 0;
parameter W42TO54 = 0;
parameter W42TO55 = 0;
parameter W42TO56 = 0;
parameter W42TO57 = 0;
parameter W42TO58 = 0;
parameter W42TO59 = 0;
parameter W42TO60 = 0;
parameter W42TO61 = 0;
parameter W42TO62 = 0;
parameter W42TO63 = 0;
parameter W42TO64 = 0;
parameter W42TO65 = 0;
parameter W42TO66 = 0;
parameter W42TO67 = 0;
parameter W42TO68 = 0;
parameter W42TO69 = 0;
parameter W42TO70 = 0;
parameter W42TO71 = 0;
parameter W42TO72 = 0;
parameter W42TO73 = 0;
parameter W42TO74 = 0;
parameter W42TO75 = 0;
parameter W42TO76 = 0;
parameter W42TO77 = 0;
parameter W42TO78 = 0;
parameter W42TO79 = 0;
parameter W42TO80 = 0;
parameter W42TO81 = 0;
parameter W42TO82 = 0;
parameter W42TO83 = 0;
parameter W42TO84 = 0;
parameter W42TO85 = 0;
parameter W42TO86 = 0;
parameter W42TO87 = 0;
parameter W42TO88 = 0;
parameter W42TO89 = 0;
parameter W42TO90 = 0;
parameter W42TO91 = 0;
parameter W42TO92 = 0;
parameter W42TO93 = 0;
parameter W42TO94 = 0;
parameter W42TO95 = 0;
parameter W42TO96 = 0;
parameter W42TO97 = 0;
parameter W42TO98 = 0;
parameter W42TO99 = 0;
parameter W43TO0 = 0;
parameter W43TO1 = 0;
parameter W43TO2 = 0;
parameter W43TO3 = 0;
parameter W43TO4 = 0;
parameter W43TO5 = 0;
parameter W43TO6 = 0;
parameter W43TO7 = 0;
parameter W43TO8 = 0;
parameter W43TO9 = 0;
parameter W43TO10 = 0;
parameter W43TO11 = 0;
parameter W43TO12 = 0;
parameter W43TO13 = 0;
parameter W43TO14 = 0;
parameter W43TO15 = 0;
parameter W43TO16 = 0;
parameter W43TO17 = 0;
parameter W43TO18 = 0;
parameter W43TO19 = 0;
parameter W43TO20 = 0;
parameter W43TO21 = 0;
parameter W43TO22 = 0;
parameter W43TO23 = 0;
parameter W43TO24 = 0;
parameter W43TO25 = 0;
parameter W43TO26 = 0;
parameter W43TO27 = 0;
parameter W43TO28 = 0;
parameter W43TO29 = 0;
parameter W43TO30 = 0;
parameter W43TO31 = 0;
parameter W43TO32 = 0;
parameter W43TO33 = 0;
parameter W43TO34 = 0;
parameter W43TO35 = 0;
parameter W43TO36 = 0;
parameter W43TO37 = 0;
parameter W43TO38 = 0;
parameter W43TO39 = 0;
parameter W43TO40 = 0;
parameter W43TO41 = 0;
parameter W43TO42 = 0;
parameter W43TO43 = 0;
parameter W43TO44 = 0;
parameter W43TO45 = 0;
parameter W43TO46 = 0;
parameter W43TO47 = 0;
parameter W43TO48 = 0;
parameter W43TO49 = 0;
parameter W43TO50 = 0;
parameter W43TO51 = 0;
parameter W43TO52 = 0;
parameter W43TO53 = 0;
parameter W43TO54 = 0;
parameter W43TO55 = 0;
parameter W43TO56 = 0;
parameter W43TO57 = 0;
parameter W43TO58 = 0;
parameter W43TO59 = 0;
parameter W43TO60 = 0;
parameter W43TO61 = 0;
parameter W43TO62 = 0;
parameter W43TO63 = 0;
parameter W43TO64 = 0;
parameter W43TO65 = 0;
parameter W43TO66 = 0;
parameter W43TO67 = 0;
parameter W43TO68 = 0;
parameter W43TO69 = 0;
parameter W43TO70 = 0;
parameter W43TO71 = 0;
parameter W43TO72 = 0;
parameter W43TO73 = 0;
parameter W43TO74 = 0;
parameter W43TO75 = 0;
parameter W43TO76 = 0;
parameter W43TO77 = 0;
parameter W43TO78 = 0;
parameter W43TO79 = 0;
parameter W43TO80 = 0;
parameter W43TO81 = 0;
parameter W43TO82 = 0;
parameter W43TO83 = 0;
parameter W43TO84 = 0;
parameter W43TO85 = 0;
parameter W43TO86 = 0;
parameter W43TO87 = 0;
parameter W43TO88 = 0;
parameter W43TO89 = 0;
parameter W43TO90 = 0;
parameter W43TO91 = 0;
parameter W43TO92 = 0;
parameter W43TO93 = 0;
parameter W43TO94 = 0;
parameter W43TO95 = 0;
parameter W43TO96 = 0;
parameter W43TO97 = 0;
parameter W43TO98 = 0;
parameter W43TO99 = 0;
parameter W44TO0 = 0;
parameter W44TO1 = 0;
parameter W44TO2 = 0;
parameter W44TO3 = 0;
parameter W44TO4 = 0;
parameter W44TO5 = 0;
parameter W44TO6 = 0;
parameter W44TO7 = 0;
parameter W44TO8 = 0;
parameter W44TO9 = 0;
parameter W44TO10 = 0;
parameter W44TO11 = 0;
parameter W44TO12 = 0;
parameter W44TO13 = 0;
parameter W44TO14 = 0;
parameter W44TO15 = 0;
parameter W44TO16 = 0;
parameter W44TO17 = 0;
parameter W44TO18 = 0;
parameter W44TO19 = 0;
parameter W44TO20 = 0;
parameter W44TO21 = 0;
parameter W44TO22 = 0;
parameter W44TO23 = 0;
parameter W44TO24 = 0;
parameter W44TO25 = 0;
parameter W44TO26 = 0;
parameter W44TO27 = 0;
parameter W44TO28 = 0;
parameter W44TO29 = 0;
parameter W44TO30 = 0;
parameter W44TO31 = 0;
parameter W44TO32 = 0;
parameter W44TO33 = 0;
parameter W44TO34 = 0;
parameter W44TO35 = 0;
parameter W44TO36 = 0;
parameter W44TO37 = 0;
parameter W44TO38 = 0;
parameter W44TO39 = 0;
parameter W44TO40 = 0;
parameter W44TO41 = 0;
parameter W44TO42 = 0;
parameter W44TO43 = 0;
parameter W44TO44 = 0;
parameter W44TO45 = 0;
parameter W44TO46 = 0;
parameter W44TO47 = 0;
parameter W44TO48 = 0;
parameter W44TO49 = 0;
parameter W44TO50 = 0;
parameter W44TO51 = 0;
parameter W44TO52 = 0;
parameter W44TO53 = 0;
parameter W44TO54 = 0;
parameter W44TO55 = 0;
parameter W44TO56 = 0;
parameter W44TO57 = 0;
parameter W44TO58 = 0;
parameter W44TO59 = 0;
parameter W44TO60 = 0;
parameter W44TO61 = 0;
parameter W44TO62 = 0;
parameter W44TO63 = 0;
parameter W44TO64 = 0;
parameter W44TO65 = 0;
parameter W44TO66 = 0;
parameter W44TO67 = 0;
parameter W44TO68 = 0;
parameter W44TO69 = 0;
parameter W44TO70 = 0;
parameter W44TO71 = 0;
parameter W44TO72 = 0;
parameter W44TO73 = 0;
parameter W44TO74 = 0;
parameter W44TO75 = 0;
parameter W44TO76 = 0;
parameter W44TO77 = 0;
parameter W44TO78 = 0;
parameter W44TO79 = 0;
parameter W44TO80 = 0;
parameter W44TO81 = 0;
parameter W44TO82 = 0;
parameter W44TO83 = 0;
parameter W44TO84 = 0;
parameter W44TO85 = 0;
parameter W44TO86 = 0;
parameter W44TO87 = 0;
parameter W44TO88 = 0;
parameter W44TO89 = 0;
parameter W44TO90 = 0;
parameter W44TO91 = 0;
parameter W44TO92 = 0;
parameter W44TO93 = 0;
parameter W44TO94 = 0;
parameter W44TO95 = 0;
parameter W44TO96 = 0;
parameter W44TO97 = 0;
parameter W44TO98 = 0;
parameter W44TO99 = 0;
parameter W45TO0 = 0;
parameter W45TO1 = 0;
parameter W45TO2 = 0;
parameter W45TO3 = 0;
parameter W45TO4 = 0;
parameter W45TO5 = 0;
parameter W45TO6 = 0;
parameter W45TO7 = 0;
parameter W45TO8 = 0;
parameter W45TO9 = 0;
parameter W45TO10 = 0;
parameter W45TO11 = 0;
parameter W45TO12 = 0;
parameter W45TO13 = 0;
parameter W45TO14 = 0;
parameter W45TO15 = 0;
parameter W45TO16 = 0;
parameter W45TO17 = 0;
parameter W45TO18 = 0;
parameter W45TO19 = 0;
parameter W45TO20 = 0;
parameter W45TO21 = 0;
parameter W45TO22 = 0;
parameter W45TO23 = 0;
parameter W45TO24 = 0;
parameter W45TO25 = 0;
parameter W45TO26 = 0;
parameter W45TO27 = 0;
parameter W45TO28 = 0;
parameter W45TO29 = 0;
parameter W45TO30 = 0;
parameter W45TO31 = 0;
parameter W45TO32 = 0;
parameter W45TO33 = 0;
parameter W45TO34 = 0;
parameter W45TO35 = 0;
parameter W45TO36 = 0;
parameter W45TO37 = 0;
parameter W45TO38 = 0;
parameter W45TO39 = 0;
parameter W45TO40 = 0;
parameter W45TO41 = 0;
parameter W45TO42 = 0;
parameter W45TO43 = 0;
parameter W45TO44 = 0;
parameter W45TO45 = 0;
parameter W45TO46 = 0;
parameter W45TO47 = 0;
parameter W45TO48 = 0;
parameter W45TO49 = 0;
parameter W45TO50 = 0;
parameter W45TO51 = 0;
parameter W45TO52 = 0;
parameter W45TO53 = 0;
parameter W45TO54 = 0;
parameter W45TO55 = 0;
parameter W45TO56 = 0;
parameter W45TO57 = 0;
parameter W45TO58 = 0;
parameter W45TO59 = 0;
parameter W45TO60 = 0;
parameter W45TO61 = 0;
parameter W45TO62 = 0;
parameter W45TO63 = 0;
parameter W45TO64 = 0;
parameter W45TO65 = 0;
parameter W45TO66 = 0;
parameter W45TO67 = 0;
parameter W45TO68 = 0;
parameter W45TO69 = 0;
parameter W45TO70 = 0;
parameter W45TO71 = 0;
parameter W45TO72 = 0;
parameter W45TO73 = 0;
parameter W45TO74 = 0;
parameter W45TO75 = 0;
parameter W45TO76 = 0;
parameter W45TO77 = 0;
parameter W45TO78 = 0;
parameter W45TO79 = 0;
parameter W45TO80 = 0;
parameter W45TO81 = 0;
parameter W45TO82 = 0;
parameter W45TO83 = 0;
parameter W45TO84 = 0;
parameter W45TO85 = 0;
parameter W45TO86 = 0;
parameter W45TO87 = 0;
parameter W45TO88 = 0;
parameter W45TO89 = 0;
parameter W45TO90 = 0;
parameter W45TO91 = 0;
parameter W45TO92 = 0;
parameter W45TO93 = 0;
parameter W45TO94 = 0;
parameter W45TO95 = 0;
parameter W45TO96 = 0;
parameter W45TO97 = 0;
parameter W45TO98 = 0;
parameter W45TO99 = 0;
parameter W46TO0 = 0;
parameter W46TO1 = 0;
parameter W46TO2 = 0;
parameter W46TO3 = 0;
parameter W46TO4 = 0;
parameter W46TO5 = 0;
parameter W46TO6 = 0;
parameter W46TO7 = 0;
parameter W46TO8 = 0;
parameter W46TO9 = 0;
parameter W46TO10 = 0;
parameter W46TO11 = 0;
parameter W46TO12 = 0;
parameter W46TO13 = 0;
parameter W46TO14 = 0;
parameter W46TO15 = 0;
parameter W46TO16 = 0;
parameter W46TO17 = 0;
parameter W46TO18 = 0;
parameter W46TO19 = 0;
parameter W46TO20 = 0;
parameter W46TO21 = 0;
parameter W46TO22 = 0;
parameter W46TO23 = 0;
parameter W46TO24 = 0;
parameter W46TO25 = 0;
parameter W46TO26 = 0;
parameter W46TO27 = 0;
parameter W46TO28 = 0;
parameter W46TO29 = 0;
parameter W46TO30 = 0;
parameter W46TO31 = 0;
parameter W46TO32 = 0;
parameter W46TO33 = 0;
parameter W46TO34 = 0;
parameter W46TO35 = 0;
parameter W46TO36 = 0;
parameter W46TO37 = 0;
parameter W46TO38 = 0;
parameter W46TO39 = 0;
parameter W46TO40 = 0;
parameter W46TO41 = 0;
parameter W46TO42 = 0;
parameter W46TO43 = 0;
parameter W46TO44 = 0;
parameter W46TO45 = 0;
parameter W46TO46 = 0;
parameter W46TO47 = 0;
parameter W46TO48 = 0;
parameter W46TO49 = 0;
parameter W46TO50 = 0;
parameter W46TO51 = 0;
parameter W46TO52 = 0;
parameter W46TO53 = 0;
parameter W46TO54 = 0;
parameter W46TO55 = 0;
parameter W46TO56 = 0;
parameter W46TO57 = 0;
parameter W46TO58 = 0;
parameter W46TO59 = 0;
parameter W46TO60 = 0;
parameter W46TO61 = 0;
parameter W46TO62 = 0;
parameter W46TO63 = 0;
parameter W46TO64 = 0;
parameter W46TO65 = 0;
parameter W46TO66 = 0;
parameter W46TO67 = 0;
parameter W46TO68 = 0;
parameter W46TO69 = 0;
parameter W46TO70 = 0;
parameter W46TO71 = 0;
parameter W46TO72 = 0;
parameter W46TO73 = 0;
parameter W46TO74 = 0;
parameter W46TO75 = 0;
parameter W46TO76 = 0;
parameter W46TO77 = 0;
parameter W46TO78 = 0;
parameter W46TO79 = 0;
parameter W46TO80 = 0;
parameter W46TO81 = 0;
parameter W46TO82 = 0;
parameter W46TO83 = 0;
parameter W46TO84 = 0;
parameter W46TO85 = 0;
parameter W46TO86 = 0;
parameter W46TO87 = 0;
parameter W46TO88 = 0;
parameter W46TO89 = 0;
parameter W46TO90 = 0;
parameter W46TO91 = 0;
parameter W46TO92 = 0;
parameter W46TO93 = 0;
parameter W46TO94 = 0;
parameter W46TO95 = 0;
parameter W46TO96 = 0;
parameter W46TO97 = 0;
parameter W46TO98 = 0;
parameter W46TO99 = 0;
parameter W47TO0 = 0;
parameter W47TO1 = 0;
parameter W47TO2 = 0;
parameter W47TO3 = 0;
parameter W47TO4 = 0;
parameter W47TO5 = 0;
parameter W47TO6 = 0;
parameter W47TO7 = 0;
parameter W47TO8 = 0;
parameter W47TO9 = 0;
parameter W47TO10 = 0;
parameter W47TO11 = 0;
parameter W47TO12 = 0;
parameter W47TO13 = 0;
parameter W47TO14 = 0;
parameter W47TO15 = 0;
parameter W47TO16 = 0;
parameter W47TO17 = 0;
parameter W47TO18 = 0;
parameter W47TO19 = 0;
parameter W47TO20 = 0;
parameter W47TO21 = 0;
parameter W47TO22 = 0;
parameter W47TO23 = 0;
parameter W47TO24 = 0;
parameter W47TO25 = 0;
parameter W47TO26 = 0;
parameter W47TO27 = 0;
parameter W47TO28 = 0;
parameter W47TO29 = 0;
parameter W47TO30 = 0;
parameter W47TO31 = 0;
parameter W47TO32 = 0;
parameter W47TO33 = 0;
parameter W47TO34 = 0;
parameter W47TO35 = 0;
parameter W47TO36 = 0;
parameter W47TO37 = 0;
parameter W47TO38 = 0;
parameter W47TO39 = 0;
parameter W47TO40 = 0;
parameter W47TO41 = 0;
parameter W47TO42 = 0;
parameter W47TO43 = 0;
parameter W47TO44 = 0;
parameter W47TO45 = 0;
parameter W47TO46 = 0;
parameter W47TO47 = 0;
parameter W47TO48 = 0;
parameter W47TO49 = 0;
parameter W47TO50 = 0;
parameter W47TO51 = 0;
parameter W47TO52 = 0;
parameter W47TO53 = 0;
parameter W47TO54 = 0;
parameter W47TO55 = 0;
parameter W47TO56 = 0;
parameter W47TO57 = 0;
parameter W47TO58 = 0;
parameter W47TO59 = 0;
parameter W47TO60 = 0;
parameter W47TO61 = 0;
parameter W47TO62 = 0;
parameter W47TO63 = 0;
parameter W47TO64 = 0;
parameter W47TO65 = 0;
parameter W47TO66 = 0;
parameter W47TO67 = 0;
parameter W47TO68 = 0;
parameter W47TO69 = 0;
parameter W47TO70 = 0;
parameter W47TO71 = 0;
parameter W47TO72 = 0;
parameter W47TO73 = 0;
parameter W47TO74 = 0;
parameter W47TO75 = 0;
parameter W47TO76 = 0;
parameter W47TO77 = 0;
parameter W47TO78 = 0;
parameter W47TO79 = 0;
parameter W47TO80 = 0;
parameter W47TO81 = 0;
parameter W47TO82 = 0;
parameter W47TO83 = 0;
parameter W47TO84 = 0;
parameter W47TO85 = 0;
parameter W47TO86 = 0;
parameter W47TO87 = 0;
parameter W47TO88 = 0;
parameter W47TO89 = 0;
parameter W47TO90 = 0;
parameter W47TO91 = 0;
parameter W47TO92 = 0;
parameter W47TO93 = 0;
parameter W47TO94 = 0;
parameter W47TO95 = 0;
parameter W47TO96 = 0;
parameter W47TO97 = 0;
parameter W47TO98 = 0;
parameter W47TO99 = 0;
parameter W48TO0 = 0;
parameter W48TO1 = 0;
parameter W48TO2 = 0;
parameter W48TO3 = 0;
parameter W48TO4 = 0;
parameter W48TO5 = 0;
parameter W48TO6 = 0;
parameter W48TO7 = 0;
parameter W48TO8 = 0;
parameter W48TO9 = 0;
parameter W48TO10 = 0;
parameter W48TO11 = 0;
parameter W48TO12 = 0;
parameter W48TO13 = 0;
parameter W48TO14 = 0;
parameter W48TO15 = 0;
parameter W48TO16 = 0;
parameter W48TO17 = 0;
parameter W48TO18 = 0;
parameter W48TO19 = 0;
parameter W48TO20 = 0;
parameter W48TO21 = 0;
parameter W48TO22 = 0;
parameter W48TO23 = 0;
parameter W48TO24 = 0;
parameter W48TO25 = 0;
parameter W48TO26 = 0;
parameter W48TO27 = 0;
parameter W48TO28 = 0;
parameter W48TO29 = 0;
parameter W48TO30 = 0;
parameter W48TO31 = 0;
parameter W48TO32 = 0;
parameter W48TO33 = 0;
parameter W48TO34 = 0;
parameter W48TO35 = 0;
parameter W48TO36 = 0;
parameter W48TO37 = 0;
parameter W48TO38 = 0;
parameter W48TO39 = 0;
parameter W48TO40 = 0;
parameter W48TO41 = 0;
parameter W48TO42 = 0;
parameter W48TO43 = 0;
parameter W48TO44 = 0;
parameter W48TO45 = 0;
parameter W48TO46 = 0;
parameter W48TO47 = 0;
parameter W48TO48 = 0;
parameter W48TO49 = 0;
parameter W48TO50 = 0;
parameter W48TO51 = 0;
parameter W48TO52 = 0;
parameter W48TO53 = 0;
parameter W48TO54 = 0;
parameter W48TO55 = 0;
parameter W48TO56 = 0;
parameter W48TO57 = 0;
parameter W48TO58 = 0;
parameter W48TO59 = 0;
parameter W48TO60 = 0;
parameter W48TO61 = 0;
parameter W48TO62 = 0;
parameter W48TO63 = 0;
parameter W48TO64 = 0;
parameter W48TO65 = 0;
parameter W48TO66 = 0;
parameter W48TO67 = 0;
parameter W48TO68 = 0;
parameter W48TO69 = 0;
parameter W48TO70 = 0;
parameter W48TO71 = 0;
parameter W48TO72 = 0;
parameter W48TO73 = 0;
parameter W48TO74 = 0;
parameter W48TO75 = 0;
parameter W48TO76 = 0;
parameter W48TO77 = 0;
parameter W48TO78 = 0;
parameter W48TO79 = 0;
parameter W48TO80 = 0;
parameter W48TO81 = 0;
parameter W48TO82 = 0;
parameter W48TO83 = 0;
parameter W48TO84 = 0;
parameter W48TO85 = 0;
parameter W48TO86 = 0;
parameter W48TO87 = 0;
parameter W48TO88 = 0;
parameter W48TO89 = 0;
parameter W48TO90 = 0;
parameter W48TO91 = 0;
parameter W48TO92 = 0;
parameter W48TO93 = 0;
parameter W48TO94 = 0;
parameter W48TO95 = 0;
parameter W48TO96 = 0;
parameter W48TO97 = 0;
parameter W48TO98 = 0;
parameter W48TO99 = 0;
parameter W49TO0 = 0;
parameter W49TO1 = 0;
parameter W49TO2 = 0;
parameter W49TO3 = 0;
parameter W49TO4 = 0;
parameter W49TO5 = 0;
parameter W49TO6 = 0;
parameter W49TO7 = 0;
parameter W49TO8 = 0;
parameter W49TO9 = 0;
parameter W49TO10 = 0;
parameter W49TO11 = 0;
parameter W49TO12 = 0;
parameter W49TO13 = 0;
parameter W49TO14 = 0;
parameter W49TO15 = 0;
parameter W49TO16 = 0;
parameter W49TO17 = 0;
parameter W49TO18 = 0;
parameter W49TO19 = 0;
parameter W49TO20 = 0;
parameter W49TO21 = 0;
parameter W49TO22 = 0;
parameter W49TO23 = 0;
parameter W49TO24 = 0;
parameter W49TO25 = 0;
parameter W49TO26 = 0;
parameter W49TO27 = 0;
parameter W49TO28 = 0;
parameter W49TO29 = 0;
parameter W49TO30 = 0;
parameter W49TO31 = 0;
parameter W49TO32 = 0;
parameter W49TO33 = 0;
parameter W49TO34 = 0;
parameter W49TO35 = 0;
parameter W49TO36 = 0;
parameter W49TO37 = 0;
parameter W49TO38 = 0;
parameter W49TO39 = 0;
parameter W49TO40 = 0;
parameter W49TO41 = 0;
parameter W49TO42 = 0;
parameter W49TO43 = 0;
parameter W49TO44 = 0;
parameter W49TO45 = 0;
parameter W49TO46 = 0;
parameter W49TO47 = 0;
parameter W49TO48 = 0;
parameter W49TO49 = 0;
parameter W49TO50 = 0;
parameter W49TO51 = 0;
parameter W49TO52 = 0;
parameter W49TO53 = 0;
parameter W49TO54 = 0;
parameter W49TO55 = 0;
parameter W49TO56 = 0;
parameter W49TO57 = 0;
parameter W49TO58 = 0;
parameter W49TO59 = 0;
parameter W49TO60 = 0;
parameter W49TO61 = 0;
parameter W49TO62 = 0;
parameter W49TO63 = 0;
parameter W49TO64 = 0;
parameter W49TO65 = 0;
parameter W49TO66 = 0;
parameter W49TO67 = 0;
parameter W49TO68 = 0;
parameter W49TO69 = 0;
parameter W49TO70 = 0;
parameter W49TO71 = 0;
parameter W49TO72 = 0;
parameter W49TO73 = 0;
parameter W49TO74 = 0;
parameter W49TO75 = 0;
parameter W49TO76 = 0;
parameter W49TO77 = 0;
parameter W49TO78 = 0;
parameter W49TO79 = 0;
parameter W49TO80 = 0;
parameter W49TO81 = 0;
parameter W49TO82 = 0;
parameter W49TO83 = 0;
parameter W49TO84 = 0;
parameter W49TO85 = 0;
parameter W49TO86 = 0;
parameter W49TO87 = 0;
parameter W49TO88 = 0;
parameter W49TO89 = 0;
parameter W49TO90 = 0;
parameter W49TO91 = 0;
parameter W49TO92 = 0;
parameter W49TO93 = 0;
parameter W49TO94 = 0;
parameter W49TO95 = 0;
parameter W49TO96 = 0;
parameter W49TO97 = 0;
parameter W49TO98 = 0;
parameter W49TO99 = 0;
parameter W50TO0 = 0;
parameter W50TO1 = 0;
parameter W50TO2 = 0;
parameter W50TO3 = 0;
parameter W50TO4 = 0;
parameter W50TO5 = 0;
parameter W50TO6 = 0;
parameter W50TO7 = 0;
parameter W50TO8 = 0;
parameter W50TO9 = 0;
parameter W50TO10 = 0;
parameter W50TO11 = 0;
parameter W50TO12 = 0;
parameter W50TO13 = 0;
parameter W50TO14 = 0;
parameter W50TO15 = 0;
parameter W50TO16 = 0;
parameter W50TO17 = 0;
parameter W50TO18 = 0;
parameter W50TO19 = 0;
parameter W50TO20 = 0;
parameter W50TO21 = 0;
parameter W50TO22 = 0;
parameter W50TO23 = 0;
parameter W50TO24 = 0;
parameter W50TO25 = 0;
parameter W50TO26 = 0;
parameter W50TO27 = 0;
parameter W50TO28 = 0;
parameter W50TO29 = 0;
parameter W50TO30 = 0;
parameter W50TO31 = 0;
parameter W50TO32 = 0;
parameter W50TO33 = 0;
parameter W50TO34 = 0;
parameter W50TO35 = 0;
parameter W50TO36 = 0;
parameter W50TO37 = 0;
parameter W50TO38 = 0;
parameter W50TO39 = 0;
parameter W50TO40 = 0;
parameter W50TO41 = 0;
parameter W50TO42 = 0;
parameter W50TO43 = 0;
parameter W50TO44 = 0;
parameter W50TO45 = 0;
parameter W50TO46 = 0;
parameter W50TO47 = 0;
parameter W50TO48 = 0;
parameter W50TO49 = 0;
parameter W50TO50 = 0;
parameter W50TO51 = 0;
parameter W50TO52 = 0;
parameter W50TO53 = 0;
parameter W50TO54 = 0;
parameter W50TO55 = 0;
parameter W50TO56 = 0;
parameter W50TO57 = 0;
parameter W50TO58 = 0;
parameter W50TO59 = 0;
parameter W50TO60 = 0;
parameter W50TO61 = 0;
parameter W50TO62 = 0;
parameter W50TO63 = 0;
parameter W50TO64 = 0;
parameter W50TO65 = 0;
parameter W50TO66 = 0;
parameter W50TO67 = 0;
parameter W50TO68 = 0;
parameter W50TO69 = 0;
parameter W50TO70 = 0;
parameter W50TO71 = 0;
parameter W50TO72 = 0;
parameter W50TO73 = 0;
parameter W50TO74 = 0;
parameter W50TO75 = 0;
parameter W50TO76 = 0;
parameter W50TO77 = 0;
parameter W50TO78 = 0;
parameter W50TO79 = 0;
parameter W50TO80 = 0;
parameter W50TO81 = 0;
parameter W50TO82 = 0;
parameter W50TO83 = 0;
parameter W50TO84 = 0;
parameter W50TO85 = 0;
parameter W50TO86 = 0;
parameter W50TO87 = 0;
parameter W50TO88 = 0;
parameter W50TO89 = 0;
parameter W50TO90 = 0;
parameter W50TO91 = 0;
parameter W50TO92 = 0;
parameter W50TO93 = 0;
parameter W50TO94 = 0;
parameter W50TO95 = 0;
parameter W50TO96 = 0;
parameter W50TO97 = 0;
parameter W50TO98 = 0;
parameter W50TO99 = 0;
parameter W51TO0 = 0;
parameter W51TO1 = 0;
parameter W51TO2 = 0;
parameter W51TO3 = 0;
parameter W51TO4 = 0;
parameter W51TO5 = 0;
parameter W51TO6 = 0;
parameter W51TO7 = 0;
parameter W51TO8 = 0;
parameter W51TO9 = 0;
parameter W51TO10 = 0;
parameter W51TO11 = 0;
parameter W51TO12 = 0;
parameter W51TO13 = 0;
parameter W51TO14 = 0;
parameter W51TO15 = 0;
parameter W51TO16 = 0;
parameter W51TO17 = 0;
parameter W51TO18 = 0;
parameter W51TO19 = 0;
parameter W51TO20 = 0;
parameter W51TO21 = 0;
parameter W51TO22 = 0;
parameter W51TO23 = 0;
parameter W51TO24 = 0;
parameter W51TO25 = 0;
parameter W51TO26 = 0;
parameter W51TO27 = 0;
parameter W51TO28 = 0;
parameter W51TO29 = 0;
parameter W51TO30 = 0;
parameter W51TO31 = 0;
parameter W51TO32 = 0;
parameter W51TO33 = 0;
parameter W51TO34 = 0;
parameter W51TO35 = 0;
parameter W51TO36 = 0;
parameter W51TO37 = 0;
parameter W51TO38 = 0;
parameter W51TO39 = 0;
parameter W51TO40 = 0;
parameter W51TO41 = 0;
parameter W51TO42 = 0;
parameter W51TO43 = 0;
parameter W51TO44 = 0;
parameter W51TO45 = 0;
parameter W51TO46 = 0;
parameter W51TO47 = 0;
parameter W51TO48 = 0;
parameter W51TO49 = 0;
parameter W51TO50 = 0;
parameter W51TO51 = 0;
parameter W51TO52 = 0;
parameter W51TO53 = 0;
parameter W51TO54 = 0;
parameter W51TO55 = 0;
parameter W51TO56 = 0;
parameter W51TO57 = 0;
parameter W51TO58 = 0;
parameter W51TO59 = 0;
parameter W51TO60 = 0;
parameter W51TO61 = 0;
parameter W51TO62 = 0;
parameter W51TO63 = 0;
parameter W51TO64 = 0;
parameter W51TO65 = 0;
parameter W51TO66 = 0;
parameter W51TO67 = 0;
parameter W51TO68 = 0;
parameter W51TO69 = 0;
parameter W51TO70 = 0;
parameter W51TO71 = 0;
parameter W51TO72 = 0;
parameter W51TO73 = 0;
parameter W51TO74 = 0;
parameter W51TO75 = 0;
parameter W51TO76 = 0;
parameter W51TO77 = 0;
parameter W51TO78 = 0;
parameter W51TO79 = 0;
parameter W51TO80 = 0;
parameter W51TO81 = 0;
parameter W51TO82 = 0;
parameter W51TO83 = 0;
parameter W51TO84 = 0;
parameter W51TO85 = 0;
parameter W51TO86 = 0;
parameter W51TO87 = 0;
parameter W51TO88 = 0;
parameter W51TO89 = 0;
parameter W51TO90 = 0;
parameter W51TO91 = 0;
parameter W51TO92 = 0;
parameter W51TO93 = 0;
parameter W51TO94 = 0;
parameter W51TO95 = 0;
parameter W51TO96 = 0;
parameter W51TO97 = 0;
parameter W51TO98 = 0;
parameter W51TO99 = 0;
parameter W52TO0 = 0;
parameter W52TO1 = 0;
parameter W52TO2 = 0;
parameter W52TO3 = 0;
parameter W52TO4 = 0;
parameter W52TO5 = 0;
parameter W52TO6 = 0;
parameter W52TO7 = 0;
parameter W52TO8 = 0;
parameter W52TO9 = 0;
parameter W52TO10 = 0;
parameter W52TO11 = 0;
parameter W52TO12 = 0;
parameter W52TO13 = 0;
parameter W52TO14 = 0;
parameter W52TO15 = 0;
parameter W52TO16 = 0;
parameter W52TO17 = 0;
parameter W52TO18 = 0;
parameter W52TO19 = 0;
parameter W52TO20 = 0;
parameter W52TO21 = 0;
parameter W52TO22 = 0;
parameter W52TO23 = 0;
parameter W52TO24 = 0;
parameter W52TO25 = 0;
parameter W52TO26 = 0;
parameter W52TO27 = 0;
parameter W52TO28 = 0;
parameter W52TO29 = 0;
parameter W52TO30 = 0;
parameter W52TO31 = 0;
parameter W52TO32 = 0;
parameter W52TO33 = 0;
parameter W52TO34 = 0;
parameter W52TO35 = 0;
parameter W52TO36 = 0;
parameter W52TO37 = 0;
parameter W52TO38 = 0;
parameter W52TO39 = 0;
parameter W52TO40 = 0;
parameter W52TO41 = 0;
parameter W52TO42 = 0;
parameter W52TO43 = 0;
parameter W52TO44 = 0;
parameter W52TO45 = 0;
parameter W52TO46 = 0;
parameter W52TO47 = 0;
parameter W52TO48 = 0;
parameter W52TO49 = 0;
parameter W52TO50 = 0;
parameter W52TO51 = 0;
parameter W52TO52 = 0;
parameter W52TO53 = 0;
parameter W52TO54 = 0;
parameter W52TO55 = 0;
parameter W52TO56 = 0;
parameter W52TO57 = 0;
parameter W52TO58 = 0;
parameter W52TO59 = 0;
parameter W52TO60 = 0;
parameter W52TO61 = 0;
parameter W52TO62 = 0;
parameter W52TO63 = 0;
parameter W52TO64 = 0;
parameter W52TO65 = 0;
parameter W52TO66 = 0;
parameter W52TO67 = 0;
parameter W52TO68 = 0;
parameter W52TO69 = 0;
parameter W52TO70 = 0;
parameter W52TO71 = 0;
parameter W52TO72 = 0;
parameter W52TO73 = 0;
parameter W52TO74 = 0;
parameter W52TO75 = 0;
parameter W52TO76 = 0;
parameter W52TO77 = 0;
parameter W52TO78 = 0;
parameter W52TO79 = 0;
parameter W52TO80 = 0;
parameter W52TO81 = 0;
parameter W52TO82 = 0;
parameter W52TO83 = 0;
parameter W52TO84 = 0;
parameter W52TO85 = 0;
parameter W52TO86 = 0;
parameter W52TO87 = 0;
parameter W52TO88 = 0;
parameter W52TO89 = 0;
parameter W52TO90 = 0;
parameter W52TO91 = 0;
parameter W52TO92 = 0;
parameter W52TO93 = 0;
parameter W52TO94 = 0;
parameter W52TO95 = 0;
parameter W52TO96 = 0;
parameter W52TO97 = 0;
parameter W52TO98 = 0;
parameter W52TO99 = 0;
parameter W53TO0 = 0;
parameter W53TO1 = 0;
parameter W53TO2 = 0;
parameter W53TO3 = 0;
parameter W53TO4 = 0;
parameter W53TO5 = 0;
parameter W53TO6 = 0;
parameter W53TO7 = 0;
parameter W53TO8 = 0;
parameter W53TO9 = 0;
parameter W53TO10 = 0;
parameter W53TO11 = 0;
parameter W53TO12 = 0;
parameter W53TO13 = 0;
parameter W53TO14 = 0;
parameter W53TO15 = 0;
parameter W53TO16 = 0;
parameter W53TO17 = 0;
parameter W53TO18 = 0;
parameter W53TO19 = 0;
parameter W53TO20 = 0;
parameter W53TO21 = 0;
parameter W53TO22 = 0;
parameter W53TO23 = 0;
parameter W53TO24 = 0;
parameter W53TO25 = 0;
parameter W53TO26 = 0;
parameter W53TO27 = 0;
parameter W53TO28 = 0;
parameter W53TO29 = 0;
parameter W53TO30 = 0;
parameter W53TO31 = 0;
parameter W53TO32 = 0;
parameter W53TO33 = 0;
parameter W53TO34 = 0;
parameter W53TO35 = 0;
parameter W53TO36 = 0;
parameter W53TO37 = 0;
parameter W53TO38 = 0;
parameter W53TO39 = 0;
parameter W53TO40 = 0;
parameter W53TO41 = 0;
parameter W53TO42 = 0;
parameter W53TO43 = 0;
parameter W53TO44 = 0;
parameter W53TO45 = 0;
parameter W53TO46 = 0;
parameter W53TO47 = 0;
parameter W53TO48 = 0;
parameter W53TO49 = 0;
parameter W53TO50 = 0;
parameter W53TO51 = 0;
parameter W53TO52 = 0;
parameter W53TO53 = 0;
parameter W53TO54 = 0;
parameter W53TO55 = 0;
parameter W53TO56 = 0;
parameter W53TO57 = 0;
parameter W53TO58 = 0;
parameter W53TO59 = 0;
parameter W53TO60 = 0;
parameter W53TO61 = 0;
parameter W53TO62 = 0;
parameter W53TO63 = 0;
parameter W53TO64 = 0;
parameter W53TO65 = 0;
parameter W53TO66 = 0;
parameter W53TO67 = 0;
parameter W53TO68 = 0;
parameter W53TO69 = 0;
parameter W53TO70 = 0;
parameter W53TO71 = 0;
parameter W53TO72 = 0;
parameter W53TO73 = 0;
parameter W53TO74 = 0;
parameter W53TO75 = 0;
parameter W53TO76 = 0;
parameter W53TO77 = 0;
parameter W53TO78 = 0;
parameter W53TO79 = 0;
parameter W53TO80 = 0;
parameter W53TO81 = 0;
parameter W53TO82 = 0;
parameter W53TO83 = 0;
parameter W53TO84 = 0;
parameter W53TO85 = 0;
parameter W53TO86 = 0;
parameter W53TO87 = 0;
parameter W53TO88 = 0;
parameter W53TO89 = 0;
parameter W53TO90 = 0;
parameter W53TO91 = 0;
parameter W53TO92 = 0;
parameter W53TO93 = 0;
parameter W53TO94 = 0;
parameter W53TO95 = 0;
parameter W53TO96 = 0;
parameter W53TO97 = 0;
parameter W53TO98 = 0;
parameter W53TO99 = 0;
parameter W54TO0 = 0;
parameter W54TO1 = 0;
parameter W54TO2 = 0;
parameter W54TO3 = 0;
parameter W54TO4 = 0;
parameter W54TO5 = 0;
parameter W54TO6 = 0;
parameter W54TO7 = 0;
parameter W54TO8 = 0;
parameter W54TO9 = 0;
parameter W54TO10 = 0;
parameter W54TO11 = 0;
parameter W54TO12 = 0;
parameter W54TO13 = 0;
parameter W54TO14 = 0;
parameter W54TO15 = 0;
parameter W54TO16 = 0;
parameter W54TO17 = 0;
parameter W54TO18 = 0;
parameter W54TO19 = 0;
parameter W54TO20 = 0;
parameter W54TO21 = 0;
parameter W54TO22 = 0;
parameter W54TO23 = 0;
parameter W54TO24 = 0;
parameter W54TO25 = 0;
parameter W54TO26 = 0;
parameter W54TO27 = 0;
parameter W54TO28 = 0;
parameter W54TO29 = 0;
parameter W54TO30 = 0;
parameter W54TO31 = 0;
parameter W54TO32 = 0;
parameter W54TO33 = 0;
parameter W54TO34 = 0;
parameter W54TO35 = 0;
parameter W54TO36 = 0;
parameter W54TO37 = 0;
parameter W54TO38 = 0;
parameter W54TO39 = 0;
parameter W54TO40 = 0;
parameter W54TO41 = 0;
parameter W54TO42 = 0;
parameter W54TO43 = 0;
parameter W54TO44 = 0;
parameter W54TO45 = 0;
parameter W54TO46 = 0;
parameter W54TO47 = 0;
parameter W54TO48 = 0;
parameter W54TO49 = 0;
parameter W54TO50 = 0;
parameter W54TO51 = 0;
parameter W54TO52 = 0;
parameter W54TO53 = 0;
parameter W54TO54 = 0;
parameter W54TO55 = 0;
parameter W54TO56 = 0;
parameter W54TO57 = 0;
parameter W54TO58 = 0;
parameter W54TO59 = 0;
parameter W54TO60 = 0;
parameter W54TO61 = 0;
parameter W54TO62 = 0;
parameter W54TO63 = 0;
parameter W54TO64 = 0;
parameter W54TO65 = 0;
parameter W54TO66 = 0;
parameter W54TO67 = 0;
parameter W54TO68 = 0;
parameter W54TO69 = 0;
parameter W54TO70 = 0;
parameter W54TO71 = 0;
parameter W54TO72 = 0;
parameter W54TO73 = 0;
parameter W54TO74 = 0;
parameter W54TO75 = 0;
parameter W54TO76 = 0;
parameter W54TO77 = 0;
parameter W54TO78 = 0;
parameter W54TO79 = 0;
parameter W54TO80 = 0;
parameter W54TO81 = 0;
parameter W54TO82 = 0;
parameter W54TO83 = 0;
parameter W54TO84 = 0;
parameter W54TO85 = 0;
parameter W54TO86 = 0;
parameter W54TO87 = 0;
parameter W54TO88 = 0;
parameter W54TO89 = 0;
parameter W54TO90 = 0;
parameter W54TO91 = 0;
parameter W54TO92 = 0;
parameter W54TO93 = 0;
parameter W54TO94 = 0;
parameter W54TO95 = 0;
parameter W54TO96 = 0;
parameter W54TO97 = 0;
parameter W54TO98 = 0;
parameter W54TO99 = 0;
parameter W55TO0 = 0;
parameter W55TO1 = 0;
parameter W55TO2 = 0;
parameter W55TO3 = 0;
parameter W55TO4 = 0;
parameter W55TO5 = 0;
parameter W55TO6 = 0;
parameter W55TO7 = 0;
parameter W55TO8 = 0;
parameter W55TO9 = 0;
parameter W55TO10 = 0;
parameter W55TO11 = 0;
parameter W55TO12 = 0;
parameter W55TO13 = 0;
parameter W55TO14 = 0;
parameter W55TO15 = 0;
parameter W55TO16 = 0;
parameter W55TO17 = 0;
parameter W55TO18 = 0;
parameter W55TO19 = 0;
parameter W55TO20 = 0;
parameter W55TO21 = 0;
parameter W55TO22 = 0;
parameter W55TO23 = 0;
parameter W55TO24 = 0;
parameter W55TO25 = 0;
parameter W55TO26 = 0;
parameter W55TO27 = 0;
parameter W55TO28 = 0;
parameter W55TO29 = 0;
parameter W55TO30 = 0;
parameter W55TO31 = 0;
parameter W55TO32 = 0;
parameter W55TO33 = 0;
parameter W55TO34 = 0;
parameter W55TO35 = 0;
parameter W55TO36 = 0;
parameter W55TO37 = 0;
parameter W55TO38 = 0;
parameter W55TO39 = 0;
parameter W55TO40 = 0;
parameter W55TO41 = 0;
parameter W55TO42 = 0;
parameter W55TO43 = 0;
parameter W55TO44 = 0;
parameter W55TO45 = 0;
parameter W55TO46 = 0;
parameter W55TO47 = 0;
parameter W55TO48 = 0;
parameter W55TO49 = 0;
parameter W55TO50 = 0;
parameter W55TO51 = 0;
parameter W55TO52 = 0;
parameter W55TO53 = 0;
parameter W55TO54 = 0;
parameter W55TO55 = 0;
parameter W55TO56 = 0;
parameter W55TO57 = 0;
parameter W55TO58 = 0;
parameter W55TO59 = 0;
parameter W55TO60 = 0;
parameter W55TO61 = 0;
parameter W55TO62 = 0;
parameter W55TO63 = 0;
parameter W55TO64 = 0;
parameter W55TO65 = 0;
parameter W55TO66 = 0;
parameter W55TO67 = 0;
parameter W55TO68 = 0;
parameter W55TO69 = 0;
parameter W55TO70 = 0;
parameter W55TO71 = 0;
parameter W55TO72 = 0;
parameter W55TO73 = 0;
parameter W55TO74 = 0;
parameter W55TO75 = 0;
parameter W55TO76 = 0;
parameter W55TO77 = 0;
parameter W55TO78 = 0;
parameter W55TO79 = 0;
parameter W55TO80 = 0;
parameter W55TO81 = 0;
parameter W55TO82 = 0;
parameter W55TO83 = 0;
parameter W55TO84 = 0;
parameter W55TO85 = 0;
parameter W55TO86 = 0;
parameter W55TO87 = 0;
parameter W55TO88 = 0;
parameter W55TO89 = 0;
parameter W55TO90 = 0;
parameter W55TO91 = 0;
parameter W55TO92 = 0;
parameter W55TO93 = 0;
parameter W55TO94 = 0;
parameter W55TO95 = 0;
parameter W55TO96 = 0;
parameter W55TO97 = 0;
parameter W55TO98 = 0;
parameter W55TO99 = 0;
parameter W56TO0 = 0;
parameter W56TO1 = 0;
parameter W56TO2 = 0;
parameter W56TO3 = 0;
parameter W56TO4 = 0;
parameter W56TO5 = 0;
parameter W56TO6 = 0;
parameter W56TO7 = 0;
parameter W56TO8 = 0;
parameter W56TO9 = 0;
parameter W56TO10 = 0;
parameter W56TO11 = 0;
parameter W56TO12 = 0;
parameter W56TO13 = 0;
parameter W56TO14 = 0;
parameter W56TO15 = 0;
parameter W56TO16 = 0;
parameter W56TO17 = 0;
parameter W56TO18 = 0;
parameter W56TO19 = 0;
parameter W56TO20 = 0;
parameter W56TO21 = 0;
parameter W56TO22 = 0;
parameter W56TO23 = 0;
parameter W56TO24 = 0;
parameter W56TO25 = 0;
parameter W56TO26 = 0;
parameter W56TO27 = 0;
parameter W56TO28 = 0;
parameter W56TO29 = 0;
parameter W56TO30 = 0;
parameter W56TO31 = 0;
parameter W56TO32 = 0;
parameter W56TO33 = 0;
parameter W56TO34 = 0;
parameter W56TO35 = 0;
parameter W56TO36 = 0;
parameter W56TO37 = 0;
parameter W56TO38 = 0;
parameter W56TO39 = 0;
parameter W56TO40 = 0;
parameter W56TO41 = 0;
parameter W56TO42 = 0;
parameter W56TO43 = 0;
parameter W56TO44 = 0;
parameter W56TO45 = 0;
parameter W56TO46 = 0;
parameter W56TO47 = 0;
parameter W56TO48 = 0;
parameter W56TO49 = 0;
parameter W56TO50 = 0;
parameter W56TO51 = 0;
parameter W56TO52 = 0;
parameter W56TO53 = 0;
parameter W56TO54 = 0;
parameter W56TO55 = 0;
parameter W56TO56 = 0;
parameter W56TO57 = 0;
parameter W56TO58 = 0;
parameter W56TO59 = 0;
parameter W56TO60 = 0;
parameter W56TO61 = 0;
parameter W56TO62 = 0;
parameter W56TO63 = 0;
parameter W56TO64 = 0;
parameter W56TO65 = 0;
parameter W56TO66 = 0;
parameter W56TO67 = 0;
parameter W56TO68 = 0;
parameter W56TO69 = 0;
parameter W56TO70 = 0;
parameter W56TO71 = 0;
parameter W56TO72 = 0;
parameter W56TO73 = 0;
parameter W56TO74 = 0;
parameter W56TO75 = 0;
parameter W56TO76 = 0;
parameter W56TO77 = 0;
parameter W56TO78 = 0;
parameter W56TO79 = 0;
parameter W56TO80 = 0;
parameter W56TO81 = 0;
parameter W56TO82 = 0;
parameter W56TO83 = 0;
parameter W56TO84 = 0;
parameter W56TO85 = 0;
parameter W56TO86 = 0;
parameter W56TO87 = 0;
parameter W56TO88 = 0;
parameter W56TO89 = 0;
parameter W56TO90 = 0;
parameter W56TO91 = 0;
parameter W56TO92 = 0;
parameter W56TO93 = 0;
parameter W56TO94 = 0;
parameter W56TO95 = 0;
parameter W56TO96 = 0;
parameter W56TO97 = 0;
parameter W56TO98 = 0;
parameter W56TO99 = 0;
parameter W57TO0 = 0;
parameter W57TO1 = 0;
parameter W57TO2 = 0;
parameter W57TO3 = 0;
parameter W57TO4 = 0;
parameter W57TO5 = 0;
parameter W57TO6 = 0;
parameter W57TO7 = 0;
parameter W57TO8 = 0;
parameter W57TO9 = 0;
parameter W57TO10 = 0;
parameter W57TO11 = 0;
parameter W57TO12 = 0;
parameter W57TO13 = 0;
parameter W57TO14 = 0;
parameter W57TO15 = 0;
parameter W57TO16 = 0;
parameter W57TO17 = 0;
parameter W57TO18 = 0;
parameter W57TO19 = 0;
parameter W57TO20 = 0;
parameter W57TO21 = 0;
parameter W57TO22 = 0;
parameter W57TO23 = 0;
parameter W57TO24 = 0;
parameter W57TO25 = 0;
parameter W57TO26 = 0;
parameter W57TO27 = 0;
parameter W57TO28 = 0;
parameter W57TO29 = 0;
parameter W57TO30 = 0;
parameter W57TO31 = 0;
parameter W57TO32 = 0;
parameter W57TO33 = 0;
parameter W57TO34 = 0;
parameter W57TO35 = 0;
parameter W57TO36 = 0;
parameter W57TO37 = 0;
parameter W57TO38 = 0;
parameter W57TO39 = 0;
parameter W57TO40 = 0;
parameter W57TO41 = 0;
parameter W57TO42 = 0;
parameter W57TO43 = 0;
parameter W57TO44 = 0;
parameter W57TO45 = 0;
parameter W57TO46 = 0;
parameter W57TO47 = 0;
parameter W57TO48 = 0;
parameter W57TO49 = 0;
parameter W57TO50 = 0;
parameter W57TO51 = 0;
parameter W57TO52 = 0;
parameter W57TO53 = 0;
parameter W57TO54 = 0;
parameter W57TO55 = 0;
parameter W57TO56 = 0;
parameter W57TO57 = 0;
parameter W57TO58 = 0;
parameter W57TO59 = 0;
parameter W57TO60 = 0;
parameter W57TO61 = 0;
parameter W57TO62 = 0;
parameter W57TO63 = 0;
parameter W57TO64 = 0;
parameter W57TO65 = 0;
parameter W57TO66 = 0;
parameter W57TO67 = 0;
parameter W57TO68 = 0;
parameter W57TO69 = 0;
parameter W57TO70 = 0;
parameter W57TO71 = 0;
parameter W57TO72 = 0;
parameter W57TO73 = 0;
parameter W57TO74 = 0;
parameter W57TO75 = 0;
parameter W57TO76 = 0;
parameter W57TO77 = 0;
parameter W57TO78 = 0;
parameter W57TO79 = 0;
parameter W57TO80 = 0;
parameter W57TO81 = 0;
parameter W57TO82 = 0;
parameter W57TO83 = 0;
parameter W57TO84 = 0;
parameter W57TO85 = 0;
parameter W57TO86 = 0;
parameter W57TO87 = 0;
parameter W57TO88 = 0;
parameter W57TO89 = 0;
parameter W57TO90 = 0;
parameter W57TO91 = 0;
parameter W57TO92 = 0;
parameter W57TO93 = 0;
parameter W57TO94 = 0;
parameter W57TO95 = 0;
parameter W57TO96 = 0;
parameter W57TO97 = 0;
parameter W57TO98 = 0;
parameter W57TO99 = 0;
parameter W58TO0 = 0;
parameter W58TO1 = 0;
parameter W58TO2 = 0;
parameter W58TO3 = 0;
parameter W58TO4 = 0;
parameter W58TO5 = 0;
parameter W58TO6 = 0;
parameter W58TO7 = 0;
parameter W58TO8 = 0;
parameter W58TO9 = 0;
parameter W58TO10 = 0;
parameter W58TO11 = 0;
parameter W58TO12 = 0;
parameter W58TO13 = 0;
parameter W58TO14 = 0;
parameter W58TO15 = 0;
parameter W58TO16 = 0;
parameter W58TO17 = 0;
parameter W58TO18 = 0;
parameter W58TO19 = 0;
parameter W58TO20 = 0;
parameter W58TO21 = 0;
parameter W58TO22 = 0;
parameter W58TO23 = 0;
parameter W58TO24 = 0;
parameter W58TO25 = 0;
parameter W58TO26 = 0;
parameter W58TO27 = 0;
parameter W58TO28 = 0;
parameter W58TO29 = 0;
parameter W58TO30 = 0;
parameter W58TO31 = 0;
parameter W58TO32 = 0;
parameter W58TO33 = 0;
parameter W58TO34 = 0;
parameter W58TO35 = 0;
parameter W58TO36 = 0;
parameter W58TO37 = 0;
parameter W58TO38 = 0;
parameter W58TO39 = 0;
parameter W58TO40 = 0;
parameter W58TO41 = 0;
parameter W58TO42 = 0;
parameter W58TO43 = 0;
parameter W58TO44 = 0;
parameter W58TO45 = 0;
parameter W58TO46 = 0;
parameter W58TO47 = 0;
parameter W58TO48 = 0;
parameter W58TO49 = 0;
parameter W58TO50 = 0;
parameter W58TO51 = 0;
parameter W58TO52 = 0;
parameter W58TO53 = 0;
parameter W58TO54 = 0;
parameter W58TO55 = 0;
parameter W58TO56 = 0;
parameter W58TO57 = 0;
parameter W58TO58 = 0;
parameter W58TO59 = 0;
parameter W58TO60 = 0;
parameter W58TO61 = 0;
parameter W58TO62 = 0;
parameter W58TO63 = 0;
parameter W58TO64 = 0;
parameter W58TO65 = 0;
parameter W58TO66 = 0;
parameter W58TO67 = 0;
parameter W58TO68 = 0;
parameter W58TO69 = 0;
parameter W58TO70 = 0;
parameter W58TO71 = 0;
parameter W58TO72 = 0;
parameter W58TO73 = 0;
parameter W58TO74 = 0;
parameter W58TO75 = 0;
parameter W58TO76 = 0;
parameter W58TO77 = 0;
parameter W58TO78 = 0;
parameter W58TO79 = 0;
parameter W58TO80 = 0;
parameter W58TO81 = 0;
parameter W58TO82 = 0;
parameter W58TO83 = 0;
parameter W58TO84 = 0;
parameter W58TO85 = 0;
parameter W58TO86 = 0;
parameter W58TO87 = 0;
parameter W58TO88 = 0;
parameter W58TO89 = 0;
parameter W58TO90 = 0;
parameter W58TO91 = 0;
parameter W58TO92 = 0;
parameter W58TO93 = 0;
parameter W58TO94 = 0;
parameter W58TO95 = 0;
parameter W58TO96 = 0;
parameter W58TO97 = 0;
parameter W58TO98 = 0;
parameter W58TO99 = 0;
parameter W59TO0 = 0;
parameter W59TO1 = 0;
parameter W59TO2 = 0;
parameter W59TO3 = 0;
parameter W59TO4 = 0;
parameter W59TO5 = 0;
parameter W59TO6 = 0;
parameter W59TO7 = 0;
parameter W59TO8 = 0;
parameter W59TO9 = 0;
parameter W59TO10 = 0;
parameter W59TO11 = 0;
parameter W59TO12 = 0;
parameter W59TO13 = 0;
parameter W59TO14 = 0;
parameter W59TO15 = 0;
parameter W59TO16 = 0;
parameter W59TO17 = 0;
parameter W59TO18 = 0;
parameter W59TO19 = 0;
parameter W59TO20 = 0;
parameter W59TO21 = 0;
parameter W59TO22 = 0;
parameter W59TO23 = 0;
parameter W59TO24 = 0;
parameter W59TO25 = 0;
parameter W59TO26 = 0;
parameter W59TO27 = 0;
parameter W59TO28 = 0;
parameter W59TO29 = 0;
parameter W59TO30 = 0;
parameter W59TO31 = 0;
parameter W59TO32 = 0;
parameter W59TO33 = 0;
parameter W59TO34 = 0;
parameter W59TO35 = 0;
parameter W59TO36 = 0;
parameter W59TO37 = 0;
parameter W59TO38 = 0;
parameter W59TO39 = 0;
parameter W59TO40 = 0;
parameter W59TO41 = 0;
parameter W59TO42 = 0;
parameter W59TO43 = 0;
parameter W59TO44 = 0;
parameter W59TO45 = 0;
parameter W59TO46 = 0;
parameter W59TO47 = 0;
parameter W59TO48 = 0;
parameter W59TO49 = 0;
parameter W59TO50 = 0;
parameter W59TO51 = 0;
parameter W59TO52 = 0;
parameter W59TO53 = 0;
parameter W59TO54 = 0;
parameter W59TO55 = 0;
parameter W59TO56 = 0;
parameter W59TO57 = 0;
parameter W59TO58 = 0;
parameter W59TO59 = 0;
parameter W59TO60 = 0;
parameter W59TO61 = 0;
parameter W59TO62 = 0;
parameter W59TO63 = 0;
parameter W59TO64 = 0;
parameter W59TO65 = 0;
parameter W59TO66 = 0;
parameter W59TO67 = 0;
parameter W59TO68 = 0;
parameter W59TO69 = 0;
parameter W59TO70 = 0;
parameter W59TO71 = 0;
parameter W59TO72 = 0;
parameter W59TO73 = 0;
parameter W59TO74 = 0;
parameter W59TO75 = 0;
parameter W59TO76 = 0;
parameter W59TO77 = 0;
parameter W59TO78 = 0;
parameter W59TO79 = 0;
parameter W59TO80 = 0;
parameter W59TO81 = 0;
parameter W59TO82 = 0;
parameter W59TO83 = 0;
parameter W59TO84 = 0;
parameter W59TO85 = 0;
parameter W59TO86 = 0;
parameter W59TO87 = 0;
parameter W59TO88 = 0;
parameter W59TO89 = 0;
parameter W59TO90 = 0;
parameter W59TO91 = 0;
parameter W59TO92 = 0;
parameter W59TO93 = 0;
parameter W59TO94 = 0;
parameter W59TO95 = 0;
parameter W59TO96 = 0;
parameter W59TO97 = 0;
parameter W59TO98 = 0;
parameter W59TO99 = 0;
parameter W60TO0 = 0;
parameter W60TO1 = 0;
parameter W60TO2 = 0;
parameter W60TO3 = 0;
parameter W60TO4 = 0;
parameter W60TO5 = 0;
parameter W60TO6 = 0;
parameter W60TO7 = 0;
parameter W60TO8 = 0;
parameter W60TO9 = 0;
parameter W60TO10 = 0;
parameter W60TO11 = 0;
parameter W60TO12 = 0;
parameter W60TO13 = 0;
parameter W60TO14 = 0;
parameter W60TO15 = 0;
parameter W60TO16 = 0;
parameter W60TO17 = 0;
parameter W60TO18 = 0;
parameter W60TO19 = 0;
parameter W60TO20 = 0;
parameter W60TO21 = 0;
parameter W60TO22 = 0;
parameter W60TO23 = 0;
parameter W60TO24 = 0;
parameter W60TO25 = 0;
parameter W60TO26 = 0;
parameter W60TO27 = 0;
parameter W60TO28 = 0;
parameter W60TO29 = 0;
parameter W60TO30 = 0;
parameter W60TO31 = 0;
parameter W60TO32 = 0;
parameter W60TO33 = 0;
parameter W60TO34 = 0;
parameter W60TO35 = 0;
parameter W60TO36 = 0;
parameter W60TO37 = 0;
parameter W60TO38 = 0;
parameter W60TO39 = 0;
parameter W60TO40 = 0;
parameter W60TO41 = 0;
parameter W60TO42 = 0;
parameter W60TO43 = 0;
parameter W60TO44 = 0;
parameter W60TO45 = 0;
parameter W60TO46 = 0;
parameter W60TO47 = 0;
parameter W60TO48 = 0;
parameter W60TO49 = 0;
parameter W60TO50 = 0;
parameter W60TO51 = 0;
parameter W60TO52 = 0;
parameter W60TO53 = 0;
parameter W60TO54 = 0;
parameter W60TO55 = 0;
parameter W60TO56 = 0;
parameter W60TO57 = 0;
parameter W60TO58 = 0;
parameter W60TO59 = 0;
parameter W60TO60 = 0;
parameter W60TO61 = 0;
parameter W60TO62 = 0;
parameter W60TO63 = 0;
parameter W60TO64 = 0;
parameter W60TO65 = 0;
parameter W60TO66 = 0;
parameter W60TO67 = 0;
parameter W60TO68 = 0;
parameter W60TO69 = 0;
parameter W60TO70 = 0;
parameter W60TO71 = 0;
parameter W60TO72 = 0;
parameter W60TO73 = 0;
parameter W60TO74 = 0;
parameter W60TO75 = 0;
parameter W60TO76 = 0;
parameter W60TO77 = 0;
parameter W60TO78 = 0;
parameter W60TO79 = 0;
parameter W60TO80 = 0;
parameter W60TO81 = 0;
parameter W60TO82 = 0;
parameter W60TO83 = 0;
parameter W60TO84 = 0;
parameter W60TO85 = 0;
parameter W60TO86 = 0;
parameter W60TO87 = 0;
parameter W60TO88 = 0;
parameter W60TO89 = 0;
parameter W60TO90 = 0;
parameter W60TO91 = 0;
parameter W60TO92 = 0;
parameter W60TO93 = 0;
parameter W60TO94 = 0;
parameter W60TO95 = 0;
parameter W60TO96 = 0;
parameter W60TO97 = 0;
parameter W60TO98 = 0;
parameter W60TO99 = 0;
parameter W61TO0 = 0;
parameter W61TO1 = 0;
parameter W61TO2 = 0;
parameter W61TO3 = 0;
parameter W61TO4 = 0;
parameter W61TO5 = 0;
parameter W61TO6 = 0;
parameter W61TO7 = 0;
parameter W61TO8 = 0;
parameter W61TO9 = 0;
parameter W61TO10 = 0;
parameter W61TO11 = 0;
parameter W61TO12 = 0;
parameter W61TO13 = 0;
parameter W61TO14 = 0;
parameter W61TO15 = 0;
parameter W61TO16 = 0;
parameter W61TO17 = 0;
parameter W61TO18 = 0;
parameter W61TO19 = 0;
parameter W61TO20 = 0;
parameter W61TO21 = 0;
parameter W61TO22 = 0;
parameter W61TO23 = 0;
parameter W61TO24 = 0;
parameter W61TO25 = 0;
parameter W61TO26 = 0;
parameter W61TO27 = 0;
parameter W61TO28 = 0;
parameter W61TO29 = 0;
parameter W61TO30 = 0;
parameter W61TO31 = 0;
parameter W61TO32 = 0;
parameter W61TO33 = 0;
parameter W61TO34 = 0;
parameter W61TO35 = 0;
parameter W61TO36 = 0;
parameter W61TO37 = 0;
parameter W61TO38 = 0;
parameter W61TO39 = 0;
parameter W61TO40 = 0;
parameter W61TO41 = 0;
parameter W61TO42 = 0;
parameter W61TO43 = 0;
parameter W61TO44 = 0;
parameter W61TO45 = 0;
parameter W61TO46 = 0;
parameter W61TO47 = 0;
parameter W61TO48 = 0;
parameter W61TO49 = 0;
parameter W61TO50 = 0;
parameter W61TO51 = 0;
parameter W61TO52 = 0;
parameter W61TO53 = 0;
parameter W61TO54 = 0;
parameter W61TO55 = 0;
parameter W61TO56 = 0;
parameter W61TO57 = 0;
parameter W61TO58 = 0;
parameter W61TO59 = 0;
parameter W61TO60 = 0;
parameter W61TO61 = 0;
parameter W61TO62 = 0;
parameter W61TO63 = 0;
parameter W61TO64 = 0;
parameter W61TO65 = 0;
parameter W61TO66 = 0;
parameter W61TO67 = 0;
parameter W61TO68 = 0;
parameter W61TO69 = 0;
parameter W61TO70 = 0;
parameter W61TO71 = 0;
parameter W61TO72 = 0;
parameter W61TO73 = 0;
parameter W61TO74 = 0;
parameter W61TO75 = 0;
parameter W61TO76 = 0;
parameter W61TO77 = 0;
parameter W61TO78 = 0;
parameter W61TO79 = 0;
parameter W61TO80 = 0;
parameter W61TO81 = 0;
parameter W61TO82 = 0;
parameter W61TO83 = 0;
parameter W61TO84 = 0;
parameter W61TO85 = 0;
parameter W61TO86 = 0;
parameter W61TO87 = 0;
parameter W61TO88 = 0;
parameter W61TO89 = 0;
parameter W61TO90 = 0;
parameter W61TO91 = 0;
parameter W61TO92 = 0;
parameter W61TO93 = 0;
parameter W61TO94 = 0;
parameter W61TO95 = 0;
parameter W61TO96 = 0;
parameter W61TO97 = 0;
parameter W61TO98 = 0;
parameter W61TO99 = 0;
parameter W62TO0 = 0;
parameter W62TO1 = 0;
parameter W62TO2 = 0;
parameter W62TO3 = 0;
parameter W62TO4 = 0;
parameter W62TO5 = 0;
parameter W62TO6 = 0;
parameter W62TO7 = 0;
parameter W62TO8 = 0;
parameter W62TO9 = 0;
parameter W62TO10 = 0;
parameter W62TO11 = 0;
parameter W62TO12 = 0;
parameter W62TO13 = 0;
parameter W62TO14 = 0;
parameter W62TO15 = 0;
parameter W62TO16 = 0;
parameter W62TO17 = 0;
parameter W62TO18 = 0;
parameter W62TO19 = 0;
parameter W62TO20 = 0;
parameter W62TO21 = 0;
parameter W62TO22 = 0;
parameter W62TO23 = 0;
parameter W62TO24 = 0;
parameter W62TO25 = 0;
parameter W62TO26 = 0;
parameter W62TO27 = 0;
parameter W62TO28 = 0;
parameter W62TO29 = 0;
parameter W62TO30 = 0;
parameter W62TO31 = 0;
parameter W62TO32 = 0;
parameter W62TO33 = 0;
parameter W62TO34 = 0;
parameter W62TO35 = 0;
parameter W62TO36 = 0;
parameter W62TO37 = 0;
parameter W62TO38 = 0;
parameter W62TO39 = 0;
parameter W62TO40 = 0;
parameter W62TO41 = 0;
parameter W62TO42 = 0;
parameter W62TO43 = 0;
parameter W62TO44 = 0;
parameter W62TO45 = 0;
parameter W62TO46 = 0;
parameter W62TO47 = 0;
parameter W62TO48 = 0;
parameter W62TO49 = 0;
parameter W62TO50 = 0;
parameter W62TO51 = 0;
parameter W62TO52 = 0;
parameter W62TO53 = 0;
parameter W62TO54 = 0;
parameter W62TO55 = 0;
parameter W62TO56 = 0;
parameter W62TO57 = 0;
parameter W62TO58 = 0;
parameter W62TO59 = 0;
parameter W62TO60 = 0;
parameter W62TO61 = 0;
parameter W62TO62 = 0;
parameter W62TO63 = 0;
parameter W62TO64 = 0;
parameter W62TO65 = 0;
parameter W62TO66 = 0;
parameter W62TO67 = 0;
parameter W62TO68 = 0;
parameter W62TO69 = 0;
parameter W62TO70 = 0;
parameter W62TO71 = 0;
parameter W62TO72 = 0;
parameter W62TO73 = 0;
parameter W62TO74 = 0;
parameter W62TO75 = 0;
parameter W62TO76 = 0;
parameter W62TO77 = 0;
parameter W62TO78 = 0;
parameter W62TO79 = 0;
parameter W62TO80 = 0;
parameter W62TO81 = 0;
parameter W62TO82 = 0;
parameter W62TO83 = 0;
parameter W62TO84 = 0;
parameter W62TO85 = 0;
parameter W62TO86 = 0;
parameter W62TO87 = 0;
parameter W62TO88 = 0;
parameter W62TO89 = 0;
parameter W62TO90 = 0;
parameter W62TO91 = 0;
parameter W62TO92 = 0;
parameter W62TO93 = 0;
parameter W62TO94 = 0;
parameter W62TO95 = 0;
parameter W62TO96 = 0;
parameter W62TO97 = 0;
parameter W62TO98 = 0;
parameter W62TO99 = 0;
parameter W63TO0 = 0;
parameter W63TO1 = 0;
parameter W63TO2 = 0;
parameter W63TO3 = 0;
parameter W63TO4 = 0;
parameter W63TO5 = 0;
parameter W63TO6 = 0;
parameter W63TO7 = 0;
parameter W63TO8 = 0;
parameter W63TO9 = 0;
parameter W63TO10 = 0;
parameter W63TO11 = 0;
parameter W63TO12 = 0;
parameter W63TO13 = 0;
parameter W63TO14 = 0;
parameter W63TO15 = 0;
parameter W63TO16 = 0;
parameter W63TO17 = 0;
parameter W63TO18 = 0;
parameter W63TO19 = 0;
parameter W63TO20 = 0;
parameter W63TO21 = 0;
parameter W63TO22 = 0;
parameter W63TO23 = 0;
parameter W63TO24 = 0;
parameter W63TO25 = 0;
parameter W63TO26 = 0;
parameter W63TO27 = 0;
parameter W63TO28 = 0;
parameter W63TO29 = 0;
parameter W63TO30 = 0;
parameter W63TO31 = 0;
parameter W63TO32 = 0;
parameter W63TO33 = 0;
parameter W63TO34 = 0;
parameter W63TO35 = 0;
parameter W63TO36 = 0;
parameter W63TO37 = 0;
parameter W63TO38 = 0;
parameter W63TO39 = 0;
parameter W63TO40 = 0;
parameter W63TO41 = 0;
parameter W63TO42 = 0;
parameter W63TO43 = 0;
parameter W63TO44 = 0;
parameter W63TO45 = 0;
parameter W63TO46 = 0;
parameter W63TO47 = 0;
parameter W63TO48 = 0;
parameter W63TO49 = 0;
parameter W63TO50 = 0;
parameter W63TO51 = 0;
parameter W63TO52 = 0;
parameter W63TO53 = 0;
parameter W63TO54 = 0;
parameter W63TO55 = 0;
parameter W63TO56 = 0;
parameter W63TO57 = 0;
parameter W63TO58 = 0;
parameter W63TO59 = 0;
parameter W63TO60 = 0;
parameter W63TO61 = 0;
parameter W63TO62 = 0;
parameter W63TO63 = 0;
parameter W63TO64 = 0;
parameter W63TO65 = 0;
parameter W63TO66 = 0;
parameter W63TO67 = 0;
parameter W63TO68 = 0;
parameter W63TO69 = 0;
parameter W63TO70 = 0;
parameter W63TO71 = 0;
parameter W63TO72 = 0;
parameter W63TO73 = 0;
parameter W63TO74 = 0;
parameter W63TO75 = 0;
parameter W63TO76 = 0;
parameter W63TO77 = 0;
parameter W63TO78 = 0;
parameter W63TO79 = 0;
parameter W63TO80 = 0;
parameter W63TO81 = 0;
parameter W63TO82 = 0;
parameter W63TO83 = 0;
parameter W63TO84 = 0;
parameter W63TO85 = 0;
parameter W63TO86 = 0;
parameter W63TO87 = 0;
parameter W63TO88 = 0;
parameter W63TO89 = 0;
parameter W63TO90 = 0;
parameter W63TO91 = 0;
parameter W63TO92 = 0;
parameter W63TO93 = 0;
parameter W63TO94 = 0;
parameter W63TO95 = 0;
parameter W63TO96 = 0;
parameter W63TO97 = 0;
parameter W63TO98 = 0;
parameter W63TO99 = 0;

input wire clk;
input wire rst;

input signed [15:0] in0;
input signed [15:0] in1;
input signed [15:0] in2;
input signed [15:0] in3;
input signed [15:0] in4;
input signed [15:0] in5;
input signed [15:0] in6;
input signed [15:0] in7;
input signed [15:0] in8;
input signed [15:0] in9;
input signed [15:0] in10;
input signed [15:0] in11;
input signed [15:0] in12;
input signed [15:0] in13;
input signed [15:0] in14;
input signed [15:0] in15;
input signed [15:0] in16;
input signed [15:0] in17;
input signed [15:0] in18;
input signed [15:0] in19;
input signed [15:0] in20;
input signed [15:0] in21;
input signed [15:0] in22;
input signed [15:0] in23;
input signed [15:0] in24;
input signed [15:0] in25;
input signed [15:0] in26;
input signed [15:0] in27;
input signed [15:0] in28;
input signed [15:0] in29;
input signed [15:0] in30;
input signed [15:0] in31;
input signed [15:0] in32;
input signed [15:0] in33;
input signed [15:0] in34;
input signed [15:0] in35;
input signed [15:0] in36;
input signed [15:0] in37;
input signed [15:0] in38;
input signed [15:0] in39;
input signed [15:0] in40;
input signed [15:0] in41;
input signed [15:0] in42;
input signed [15:0] in43;
input signed [15:0] in44;
input signed [15:0] in45;
input signed [15:0] in46;
input signed [15:0] in47;
input signed [15:0] in48;
input signed [15:0] in49;
input signed [15:0] in50;
input signed [15:0] in51;
input signed [15:0] in52;
input signed [15:0] in53;
input signed [15:0] in54;
input signed [15:0] in55;
input signed [15:0] in56;
input signed [15:0] in57;
input signed [15:0] in58;
input signed [15:0] in59;
input signed [15:0] in60;
input signed [15:0] in61;
input signed [15:0] in62;
input signed [15:0] in63;

output signed [15:0] out0;
output signed [15:0] out1;
output signed [15:0] out2;
output signed [15:0] out3;
output signed [15:0] out4;
output signed [15:0] out5;
output signed [15:0] out6;
output signed [15:0] out7;
output signed [15:0] out8;
output signed [15:0] out9;
output signed [15:0] out10;
output signed [15:0] out11;
output signed [15:0] out12;
output signed [15:0] out13;
output signed [15:0] out14;
output signed [15:0] out15;
output signed [15:0] out16;
output signed [15:0] out17;
output signed [15:0] out18;
output signed [15:0] out19;
output signed [15:0] out20;
output signed [15:0] out21;
output signed [15:0] out22;
output signed [15:0] out23;
output signed [15:0] out24;
output signed [15:0] out25;
output signed [15:0] out26;
output signed [15:0] out27;
output signed [15:0] out28;
output signed [15:0] out29;
output signed [15:0] out30;
output signed [15:0] out31;
output signed [15:0] out32;
output signed [15:0] out33;
output signed [15:0] out34;
output signed [15:0] out35;
output signed [15:0] out36;
output signed [15:0] out37;
output signed [15:0] out38;
output signed [15:0] out39;
output signed [15:0] out40;
output signed [15:0] out41;
output signed [15:0] out42;
output signed [15:0] out43;
output signed [15:0] out44;
output signed [15:0] out45;
output signed [15:0] out46;
output signed [15:0] out47;
output signed [15:0] out48;
output signed [15:0] out49;
output signed [15:0] out50;
output signed [15:0] out51;
output signed [15:0] out52;
output signed [15:0] out53;
output signed [15:0] out54;
output signed [15:0] out55;
output signed [15:0] out56;
output signed [15:0] out57;
output signed [15:0] out58;
output signed [15:0] out59;
output signed [15:0] out60;
output signed [15:0] out61;
output signed [15:0] out62;
output signed [15:0] out63;
output signed [15:0] out64;
output signed [15:0] out65;
output signed [15:0] out66;
output signed [15:0] out67;
output signed [15:0] out68;
output signed [15:0] out69;
output signed [15:0] out70;
output signed [15:0] out71;
output signed [15:0] out72;
output signed [15:0] out73;
output signed [15:0] out74;
output signed [15:0] out75;
output signed [15:0] out76;
output signed [15:0] out77;
output signed [15:0] out78;
output signed [15:0] out79;
output signed [15:0] out80;
output signed [15:0] out81;
output signed [15:0] out82;
output signed [15:0] out83;
output signed [15:0] out84;
output signed [15:0] out85;
output signed [15:0] out86;
output signed [15:0] out87;
output signed [15:0] out88;
output signed [15:0] out89;
output signed [15:0] out90;
output signed [15:0] out91;
output signed [15:0] out92;
output signed [15:0] out93;
output signed [15:0] out94;
output signed [15:0] out95;
output signed [15:0] out96;
output signed [15:0] out97;
output signed [15:0] out98;
output signed [15:0] out99;

neuron64in #(.W0(W0TO0), .W1(W1TO0), .W2(W2TO0), .W3(W3TO0), .W4(W4TO0), .W5(W5TO0), .W6(W6TO0), .W7(W7TO0), .W8(W8TO0), .W9(W9TO0), .W10(W10TO0), .W11(W11TO0), .W12(W12TO0), .W13(W13TO0), .W14(W14TO0), .W15(W15TO0), .W16(W16TO0), .W17(W17TO0), .W18(W18TO0), .W19(W19TO0), .W20(W20TO0), .W21(W21TO0), .W22(W22TO0), .W23(W23TO0), .W24(W24TO0), .W25(W25TO0), .W26(W26TO0), .W27(W27TO0), .W28(W28TO0), .W29(W29TO0), .W30(W30TO0), .W31(W31TO0), .W32(W32TO0), .W33(W33TO0), .W34(W34TO0), .W35(W35TO0), .W36(W36TO0), .W37(W37TO0), .W38(W38TO0), .W39(W39TO0), .W40(W40TO0), .W41(W41TO0), .W42(W42TO0), .W43(W43TO0), .W44(W44TO0), .W45(W45TO0), .W46(W46TO0), .W47(W47TO0), .W48(W48TO0), .W49(W49TO0), .W50(W50TO0), .W51(W51TO0), .W52(W52TO0), .W53(W53TO0), .W54(W54TO0), .W55(W55TO0), .W56(W56TO0), .W57(W57TO0), .W58(W58TO0), .W59(W59TO0), .W60(W60TO0), .W61(W61TO0), .W62(W62TO0), .W63(W63TO0)) neuron0(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out0));
neuron64in #(.W0(W0TO1), .W1(W1TO1), .W2(W2TO1), .W3(W3TO1), .W4(W4TO1), .W5(W5TO1), .W6(W6TO1), .W7(W7TO1), .W8(W8TO1), .W9(W9TO1), .W10(W10TO1), .W11(W11TO1), .W12(W12TO1), .W13(W13TO1), .W14(W14TO1), .W15(W15TO1), .W16(W16TO1), .W17(W17TO1), .W18(W18TO1), .W19(W19TO1), .W20(W20TO1), .W21(W21TO1), .W22(W22TO1), .W23(W23TO1), .W24(W24TO1), .W25(W25TO1), .W26(W26TO1), .W27(W27TO1), .W28(W28TO1), .W29(W29TO1), .W30(W30TO1), .W31(W31TO1), .W32(W32TO1), .W33(W33TO1), .W34(W34TO1), .W35(W35TO1), .W36(W36TO1), .W37(W37TO1), .W38(W38TO1), .W39(W39TO1), .W40(W40TO1), .W41(W41TO1), .W42(W42TO1), .W43(W43TO1), .W44(W44TO1), .W45(W45TO1), .W46(W46TO1), .W47(W47TO1), .W48(W48TO1), .W49(W49TO1), .W50(W50TO1), .W51(W51TO1), .W52(W52TO1), .W53(W53TO1), .W54(W54TO1), .W55(W55TO1), .W56(W56TO1), .W57(W57TO1), .W58(W58TO1), .W59(W59TO1), .W60(W60TO1), .W61(W61TO1), .W62(W62TO1), .W63(W63TO1)) neuron1(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out1));
neuron64in #(.W0(W0TO2), .W1(W1TO2), .W2(W2TO2), .W3(W3TO2), .W4(W4TO2), .W5(W5TO2), .W6(W6TO2), .W7(W7TO2), .W8(W8TO2), .W9(W9TO2), .W10(W10TO2), .W11(W11TO2), .W12(W12TO2), .W13(W13TO2), .W14(W14TO2), .W15(W15TO2), .W16(W16TO2), .W17(W17TO2), .W18(W18TO2), .W19(W19TO2), .W20(W20TO2), .W21(W21TO2), .W22(W22TO2), .W23(W23TO2), .W24(W24TO2), .W25(W25TO2), .W26(W26TO2), .W27(W27TO2), .W28(W28TO2), .W29(W29TO2), .W30(W30TO2), .W31(W31TO2), .W32(W32TO2), .W33(W33TO2), .W34(W34TO2), .W35(W35TO2), .W36(W36TO2), .W37(W37TO2), .W38(W38TO2), .W39(W39TO2), .W40(W40TO2), .W41(W41TO2), .W42(W42TO2), .W43(W43TO2), .W44(W44TO2), .W45(W45TO2), .W46(W46TO2), .W47(W47TO2), .W48(W48TO2), .W49(W49TO2), .W50(W50TO2), .W51(W51TO2), .W52(W52TO2), .W53(W53TO2), .W54(W54TO2), .W55(W55TO2), .W56(W56TO2), .W57(W57TO2), .W58(W58TO2), .W59(W59TO2), .W60(W60TO2), .W61(W61TO2), .W62(W62TO2), .W63(W63TO2)) neuron2(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out2));
neuron64in #(.W0(W0TO3), .W1(W1TO3), .W2(W2TO3), .W3(W3TO3), .W4(W4TO3), .W5(W5TO3), .W6(W6TO3), .W7(W7TO3), .W8(W8TO3), .W9(W9TO3), .W10(W10TO3), .W11(W11TO3), .W12(W12TO3), .W13(W13TO3), .W14(W14TO3), .W15(W15TO3), .W16(W16TO3), .W17(W17TO3), .W18(W18TO3), .W19(W19TO3), .W20(W20TO3), .W21(W21TO3), .W22(W22TO3), .W23(W23TO3), .W24(W24TO3), .W25(W25TO3), .W26(W26TO3), .W27(W27TO3), .W28(W28TO3), .W29(W29TO3), .W30(W30TO3), .W31(W31TO3), .W32(W32TO3), .W33(W33TO3), .W34(W34TO3), .W35(W35TO3), .W36(W36TO3), .W37(W37TO3), .W38(W38TO3), .W39(W39TO3), .W40(W40TO3), .W41(W41TO3), .W42(W42TO3), .W43(W43TO3), .W44(W44TO3), .W45(W45TO3), .W46(W46TO3), .W47(W47TO3), .W48(W48TO3), .W49(W49TO3), .W50(W50TO3), .W51(W51TO3), .W52(W52TO3), .W53(W53TO3), .W54(W54TO3), .W55(W55TO3), .W56(W56TO3), .W57(W57TO3), .W58(W58TO3), .W59(W59TO3), .W60(W60TO3), .W61(W61TO3), .W62(W62TO3), .W63(W63TO3)) neuron3(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out3));
neuron64in #(.W0(W0TO4), .W1(W1TO4), .W2(W2TO4), .W3(W3TO4), .W4(W4TO4), .W5(W5TO4), .W6(W6TO4), .W7(W7TO4), .W8(W8TO4), .W9(W9TO4), .W10(W10TO4), .W11(W11TO4), .W12(W12TO4), .W13(W13TO4), .W14(W14TO4), .W15(W15TO4), .W16(W16TO4), .W17(W17TO4), .W18(W18TO4), .W19(W19TO4), .W20(W20TO4), .W21(W21TO4), .W22(W22TO4), .W23(W23TO4), .W24(W24TO4), .W25(W25TO4), .W26(W26TO4), .W27(W27TO4), .W28(W28TO4), .W29(W29TO4), .W30(W30TO4), .W31(W31TO4), .W32(W32TO4), .W33(W33TO4), .W34(W34TO4), .W35(W35TO4), .W36(W36TO4), .W37(W37TO4), .W38(W38TO4), .W39(W39TO4), .W40(W40TO4), .W41(W41TO4), .W42(W42TO4), .W43(W43TO4), .W44(W44TO4), .W45(W45TO4), .W46(W46TO4), .W47(W47TO4), .W48(W48TO4), .W49(W49TO4), .W50(W50TO4), .W51(W51TO4), .W52(W52TO4), .W53(W53TO4), .W54(W54TO4), .W55(W55TO4), .W56(W56TO4), .W57(W57TO4), .W58(W58TO4), .W59(W59TO4), .W60(W60TO4), .W61(W61TO4), .W62(W62TO4), .W63(W63TO4)) neuron4(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out4));
neuron64in #(.W0(W0TO5), .W1(W1TO5), .W2(W2TO5), .W3(W3TO5), .W4(W4TO5), .W5(W5TO5), .W6(W6TO5), .W7(W7TO5), .W8(W8TO5), .W9(W9TO5), .W10(W10TO5), .W11(W11TO5), .W12(W12TO5), .W13(W13TO5), .W14(W14TO5), .W15(W15TO5), .W16(W16TO5), .W17(W17TO5), .W18(W18TO5), .W19(W19TO5), .W20(W20TO5), .W21(W21TO5), .W22(W22TO5), .W23(W23TO5), .W24(W24TO5), .W25(W25TO5), .W26(W26TO5), .W27(W27TO5), .W28(W28TO5), .W29(W29TO5), .W30(W30TO5), .W31(W31TO5), .W32(W32TO5), .W33(W33TO5), .W34(W34TO5), .W35(W35TO5), .W36(W36TO5), .W37(W37TO5), .W38(W38TO5), .W39(W39TO5), .W40(W40TO5), .W41(W41TO5), .W42(W42TO5), .W43(W43TO5), .W44(W44TO5), .W45(W45TO5), .W46(W46TO5), .W47(W47TO5), .W48(W48TO5), .W49(W49TO5), .W50(W50TO5), .W51(W51TO5), .W52(W52TO5), .W53(W53TO5), .W54(W54TO5), .W55(W55TO5), .W56(W56TO5), .W57(W57TO5), .W58(W58TO5), .W59(W59TO5), .W60(W60TO5), .W61(W61TO5), .W62(W62TO5), .W63(W63TO5)) neuron5(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out5));
neuron64in #(.W0(W0TO6), .W1(W1TO6), .W2(W2TO6), .W3(W3TO6), .W4(W4TO6), .W5(W5TO6), .W6(W6TO6), .W7(W7TO6), .W8(W8TO6), .W9(W9TO6), .W10(W10TO6), .W11(W11TO6), .W12(W12TO6), .W13(W13TO6), .W14(W14TO6), .W15(W15TO6), .W16(W16TO6), .W17(W17TO6), .W18(W18TO6), .W19(W19TO6), .W20(W20TO6), .W21(W21TO6), .W22(W22TO6), .W23(W23TO6), .W24(W24TO6), .W25(W25TO6), .W26(W26TO6), .W27(W27TO6), .W28(W28TO6), .W29(W29TO6), .W30(W30TO6), .W31(W31TO6), .W32(W32TO6), .W33(W33TO6), .W34(W34TO6), .W35(W35TO6), .W36(W36TO6), .W37(W37TO6), .W38(W38TO6), .W39(W39TO6), .W40(W40TO6), .W41(W41TO6), .W42(W42TO6), .W43(W43TO6), .W44(W44TO6), .W45(W45TO6), .W46(W46TO6), .W47(W47TO6), .W48(W48TO6), .W49(W49TO6), .W50(W50TO6), .W51(W51TO6), .W52(W52TO6), .W53(W53TO6), .W54(W54TO6), .W55(W55TO6), .W56(W56TO6), .W57(W57TO6), .W58(W58TO6), .W59(W59TO6), .W60(W60TO6), .W61(W61TO6), .W62(W62TO6), .W63(W63TO6)) neuron6(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out6));
neuron64in #(.W0(W0TO7), .W1(W1TO7), .W2(W2TO7), .W3(W3TO7), .W4(W4TO7), .W5(W5TO7), .W6(W6TO7), .W7(W7TO7), .W8(W8TO7), .W9(W9TO7), .W10(W10TO7), .W11(W11TO7), .W12(W12TO7), .W13(W13TO7), .W14(W14TO7), .W15(W15TO7), .W16(W16TO7), .W17(W17TO7), .W18(W18TO7), .W19(W19TO7), .W20(W20TO7), .W21(W21TO7), .W22(W22TO7), .W23(W23TO7), .W24(W24TO7), .W25(W25TO7), .W26(W26TO7), .W27(W27TO7), .W28(W28TO7), .W29(W29TO7), .W30(W30TO7), .W31(W31TO7), .W32(W32TO7), .W33(W33TO7), .W34(W34TO7), .W35(W35TO7), .W36(W36TO7), .W37(W37TO7), .W38(W38TO7), .W39(W39TO7), .W40(W40TO7), .W41(W41TO7), .W42(W42TO7), .W43(W43TO7), .W44(W44TO7), .W45(W45TO7), .W46(W46TO7), .W47(W47TO7), .W48(W48TO7), .W49(W49TO7), .W50(W50TO7), .W51(W51TO7), .W52(W52TO7), .W53(W53TO7), .W54(W54TO7), .W55(W55TO7), .W56(W56TO7), .W57(W57TO7), .W58(W58TO7), .W59(W59TO7), .W60(W60TO7), .W61(W61TO7), .W62(W62TO7), .W63(W63TO7)) neuron7(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out7));
neuron64in #(.W0(W0TO8), .W1(W1TO8), .W2(W2TO8), .W3(W3TO8), .W4(W4TO8), .W5(W5TO8), .W6(W6TO8), .W7(W7TO8), .W8(W8TO8), .W9(W9TO8), .W10(W10TO8), .W11(W11TO8), .W12(W12TO8), .W13(W13TO8), .W14(W14TO8), .W15(W15TO8), .W16(W16TO8), .W17(W17TO8), .W18(W18TO8), .W19(W19TO8), .W20(W20TO8), .W21(W21TO8), .W22(W22TO8), .W23(W23TO8), .W24(W24TO8), .W25(W25TO8), .W26(W26TO8), .W27(W27TO8), .W28(W28TO8), .W29(W29TO8), .W30(W30TO8), .W31(W31TO8), .W32(W32TO8), .W33(W33TO8), .W34(W34TO8), .W35(W35TO8), .W36(W36TO8), .W37(W37TO8), .W38(W38TO8), .W39(W39TO8), .W40(W40TO8), .W41(W41TO8), .W42(W42TO8), .W43(W43TO8), .W44(W44TO8), .W45(W45TO8), .W46(W46TO8), .W47(W47TO8), .W48(W48TO8), .W49(W49TO8), .W50(W50TO8), .W51(W51TO8), .W52(W52TO8), .W53(W53TO8), .W54(W54TO8), .W55(W55TO8), .W56(W56TO8), .W57(W57TO8), .W58(W58TO8), .W59(W59TO8), .W60(W60TO8), .W61(W61TO8), .W62(W62TO8), .W63(W63TO8)) neuron8(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out8));
neuron64in #(.W0(W0TO9), .W1(W1TO9), .W2(W2TO9), .W3(W3TO9), .W4(W4TO9), .W5(W5TO9), .W6(W6TO9), .W7(W7TO9), .W8(W8TO9), .W9(W9TO9), .W10(W10TO9), .W11(W11TO9), .W12(W12TO9), .W13(W13TO9), .W14(W14TO9), .W15(W15TO9), .W16(W16TO9), .W17(W17TO9), .W18(W18TO9), .W19(W19TO9), .W20(W20TO9), .W21(W21TO9), .W22(W22TO9), .W23(W23TO9), .W24(W24TO9), .W25(W25TO9), .W26(W26TO9), .W27(W27TO9), .W28(W28TO9), .W29(W29TO9), .W30(W30TO9), .W31(W31TO9), .W32(W32TO9), .W33(W33TO9), .W34(W34TO9), .W35(W35TO9), .W36(W36TO9), .W37(W37TO9), .W38(W38TO9), .W39(W39TO9), .W40(W40TO9), .W41(W41TO9), .W42(W42TO9), .W43(W43TO9), .W44(W44TO9), .W45(W45TO9), .W46(W46TO9), .W47(W47TO9), .W48(W48TO9), .W49(W49TO9), .W50(W50TO9), .W51(W51TO9), .W52(W52TO9), .W53(W53TO9), .W54(W54TO9), .W55(W55TO9), .W56(W56TO9), .W57(W57TO9), .W58(W58TO9), .W59(W59TO9), .W60(W60TO9), .W61(W61TO9), .W62(W62TO9), .W63(W63TO9)) neuron9(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out9));
neuron64in #(.W0(W0TO10), .W1(W1TO10), .W2(W2TO10), .W3(W3TO10), .W4(W4TO10), .W5(W5TO10), .W6(W6TO10), .W7(W7TO10), .W8(W8TO10), .W9(W9TO10), .W10(W10TO10), .W11(W11TO10), .W12(W12TO10), .W13(W13TO10), .W14(W14TO10), .W15(W15TO10), .W16(W16TO10), .W17(W17TO10), .W18(W18TO10), .W19(W19TO10), .W20(W20TO10), .W21(W21TO10), .W22(W22TO10), .W23(W23TO10), .W24(W24TO10), .W25(W25TO10), .W26(W26TO10), .W27(W27TO10), .W28(W28TO10), .W29(W29TO10), .W30(W30TO10), .W31(W31TO10), .W32(W32TO10), .W33(W33TO10), .W34(W34TO10), .W35(W35TO10), .W36(W36TO10), .W37(W37TO10), .W38(W38TO10), .W39(W39TO10), .W40(W40TO10), .W41(W41TO10), .W42(W42TO10), .W43(W43TO10), .W44(W44TO10), .W45(W45TO10), .W46(W46TO10), .W47(W47TO10), .W48(W48TO10), .W49(W49TO10), .W50(W50TO10), .W51(W51TO10), .W52(W52TO10), .W53(W53TO10), .W54(W54TO10), .W55(W55TO10), .W56(W56TO10), .W57(W57TO10), .W58(W58TO10), .W59(W59TO10), .W60(W60TO10), .W61(W61TO10), .W62(W62TO10), .W63(W63TO10)) neuron10(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out10));
neuron64in #(.W0(W0TO11), .W1(W1TO11), .W2(W2TO11), .W3(W3TO11), .W4(W4TO11), .W5(W5TO11), .W6(W6TO11), .W7(W7TO11), .W8(W8TO11), .W9(W9TO11), .W10(W10TO11), .W11(W11TO11), .W12(W12TO11), .W13(W13TO11), .W14(W14TO11), .W15(W15TO11), .W16(W16TO11), .W17(W17TO11), .W18(W18TO11), .W19(W19TO11), .W20(W20TO11), .W21(W21TO11), .W22(W22TO11), .W23(W23TO11), .W24(W24TO11), .W25(W25TO11), .W26(W26TO11), .W27(W27TO11), .W28(W28TO11), .W29(W29TO11), .W30(W30TO11), .W31(W31TO11), .W32(W32TO11), .W33(W33TO11), .W34(W34TO11), .W35(W35TO11), .W36(W36TO11), .W37(W37TO11), .W38(W38TO11), .W39(W39TO11), .W40(W40TO11), .W41(W41TO11), .W42(W42TO11), .W43(W43TO11), .W44(W44TO11), .W45(W45TO11), .W46(W46TO11), .W47(W47TO11), .W48(W48TO11), .W49(W49TO11), .W50(W50TO11), .W51(W51TO11), .W52(W52TO11), .W53(W53TO11), .W54(W54TO11), .W55(W55TO11), .W56(W56TO11), .W57(W57TO11), .W58(W58TO11), .W59(W59TO11), .W60(W60TO11), .W61(W61TO11), .W62(W62TO11), .W63(W63TO11)) neuron11(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out11));
neuron64in #(.W0(W0TO12), .W1(W1TO12), .W2(W2TO12), .W3(W3TO12), .W4(W4TO12), .W5(W5TO12), .W6(W6TO12), .W7(W7TO12), .W8(W8TO12), .W9(W9TO12), .W10(W10TO12), .W11(W11TO12), .W12(W12TO12), .W13(W13TO12), .W14(W14TO12), .W15(W15TO12), .W16(W16TO12), .W17(W17TO12), .W18(W18TO12), .W19(W19TO12), .W20(W20TO12), .W21(W21TO12), .W22(W22TO12), .W23(W23TO12), .W24(W24TO12), .W25(W25TO12), .W26(W26TO12), .W27(W27TO12), .W28(W28TO12), .W29(W29TO12), .W30(W30TO12), .W31(W31TO12), .W32(W32TO12), .W33(W33TO12), .W34(W34TO12), .W35(W35TO12), .W36(W36TO12), .W37(W37TO12), .W38(W38TO12), .W39(W39TO12), .W40(W40TO12), .W41(W41TO12), .W42(W42TO12), .W43(W43TO12), .W44(W44TO12), .W45(W45TO12), .W46(W46TO12), .W47(W47TO12), .W48(W48TO12), .W49(W49TO12), .W50(W50TO12), .W51(W51TO12), .W52(W52TO12), .W53(W53TO12), .W54(W54TO12), .W55(W55TO12), .W56(W56TO12), .W57(W57TO12), .W58(W58TO12), .W59(W59TO12), .W60(W60TO12), .W61(W61TO12), .W62(W62TO12), .W63(W63TO12)) neuron12(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out12));
neuron64in #(.W0(W0TO13), .W1(W1TO13), .W2(W2TO13), .W3(W3TO13), .W4(W4TO13), .W5(W5TO13), .W6(W6TO13), .W7(W7TO13), .W8(W8TO13), .W9(W9TO13), .W10(W10TO13), .W11(W11TO13), .W12(W12TO13), .W13(W13TO13), .W14(W14TO13), .W15(W15TO13), .W16(W16TO13), .W17(W17TO13), .W18(W18TO13), .W19(W19TO13), .W20(W20TO13), .W21(W21TO13), .W22(W22TO13), .W23(W23TO13), .W24(W24TO13), .W25(W25TO13), .W26(W26TO13), .W27(W27TO13), .W28(W28TO13), .W29(W29TO13), .W30(W30TO13), .W31(W31TO13), .W32(W32TO13), .W33(W33TO13), .W34(W34TO13), .W35(W35TO13), .W36(W36TO13), .W37(W37TO13), .W38(W38TO13), .W39(W39TO13), .W40(W40TO13), .W41(W41TO13), .W42(W42TO13), .W43(W43TO13), .W44(W44TO13), .W45(W45TO13), .W46(W46TO13), .W47(W47TO13), .W48(W48TO13), .W49(W49TO13), .W50(W50TO13), .W51(W51TO13), .W52(W52TO13), .W53(W53TO13), .W54(W54TO13), .W55(W55TO13), .W56(W56TO13), .W57(W57TO13), .W58(W58TO13), .W59(W59TO13), .W60(W60TO13), .W61(W61TO13), .W62(W62TO13), .W63(W63TO13)) neuron13(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out13));
neuron64in #(.W0(W0TO14), .W1(W1TO14), .W2(W2TO14), .W3(W3TO14), .W4(W4TO14), .W5(W5TO14), .W6(W6TO14), .W7(W7TO14), .W8(W8TO14), .W9(W9TO14), .W10(W10TO14), .W11(W11TO14), .W12(W12TO14), .W13(W13TO14), .W14(W14TO14), .W15(W15TO14), .W16(W16TO14), .W17(W17TO14), .W18(W18TO14), .W19(W19TO14), .W20(W20TO14), .W21(W21TO14), .W22(W22TO14), .W23(W23TO14), .W24(W24TO14), .W25(W25TO14), .W26(W26TO14), .W27(W27TO14), .W28(W28TO14), .W29(W29TO14), .W30(W30TO14), .W31(W31TO14), .W32(W32TO14), .W33(W33TO14), .W34(W34TO14), .W35(W35TO14), .W36(W36TO14), .W37(W37TO14), .W38(W38TO14), .W39(W39TO14), .W40(W40TO14), .W41(W41TO14), .W42(W42TO14), .W43(W43TO14), .W44(W44TO14), .W45(W45TO14), .W46(W46TO14), .W47(W47TO14), .W48(W48TO14), .W49(W49TO14), .W50(W50TO14), .W51(W51TO14), .W52(W52TO14), .W53(W53TO14), .W54(W54TO14), .W55(W55TO14), .W56(W56TO14), .W57(W57TO14), .W58(W58TO14), .W59(W59TO14), .W60(W60TO14), .W61(W61TO14), .W62(W62TO14), .W63(W63TO14)) neuron14(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out14));
neuron64in #(.W0(W0TO15), .W1(W1TO15), .W2(W2TO15), .W3(W3TO15), .W4(W4TO15), .W5(W5TO15), .W6(W6TO15), .W7(W7TO15), .W8(W8TO15), .W9(W9TO15), .W10(W10TO15), .W11(W11TO15), .W12(W12TO15), .W13(W13TO15), .W14(W14TO15), .W15(W15TO15), .W16(W16TO15), .W17(W17TO15), .W18(W18TO15), .W19(W19TO15), .W20(W20TO15), .W21(W21TO15), .W22(W22TO15), .W23(W23TO15), .W24(W24TO15), .W25(W25TO15), .W26(W26TO15), .W27(W27TO15), .W28(W28TO15), .W29(W29TO15), .W30(W30TO15), .W31(W31TO15), .W32(W32TO15), .W33(W33TO15), .W34(W34TO15), .W35(W35TO15), .W36(W36TO15), .W37(W37TO15), .W38(W38TO15), .W39(W39TO15), .W40(W40TO15), .W41(W41TO15), .W42(W42TO15), .W43(W43TO15), .W44(W44TO15), .W45(W45TO15), .W46(W46TO15), .W47(W47TO15), .W48(W48TO15), .W49(W49TO15), .W50(W50TO15), .W51(W51TO15), .W52(W52TO15), .W53(W53TO15), .W54(W54TO15), .W55(W55TO15), .W56(W56TO15), .W57(W57TO15), .W58(W58TO15), .W59(W59TO15), .W60(W60TO15), .W61(W61TO15), .W62(W62TO15), .W63(W63TO15)) neuron15(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out15));
neuron64in #(.W0(W0TO16), .W1(W1TO16), .W2(W2TO16), .W3(W3TO16), .W4(W4TO16), .W5(W5TO16), .W6(W6TO16), .W7(W7TO16), .W8(W8TO16), .W9(W9TO16), .W10(W10TO16), .W11(W11TO16), .W12(W12TO16), .W13(W13TO16), .W14(W14TO16), .W15(W15TO16), .W16(W16TO16), .W17(W17TO16), .W18(W18TO16), .W19(W19TO16), .W20(W20TO16), .W21(W21TO16), .W22(W22TO16), .W23(W23TO16), .W24(W24TO16), .W25(W25TO16), .W26(W26TO16), .W27(W27TO16), .W28(W28TO16), .W29(W29TO16), .W30(W30TO16), .W31(W31TO16), .W32(W32TO16), .W33(W33TO16), .W34(W34TO16), .W35(W35TO16), .W36(W36TO16), .W37(W37TO16), .W38(W38TO16), .W39(W39TO16), .W40(W40TO16), .W41(W41TO16), .W42(W42TO16), .W43(W43TO16), .W44(W44TO16), .W45(W45TO16), .W46(W46TO16), .W47(W47TO16), .W48(W48TO16), .W49(W49TO16), .W50(W50TO16), .W51(W51TO16), .W52(W52TO16), .W53(W53TO16), .W54(W54TO16), .W55(W55TO16), .W56(W56TO16), .W57(W57TO16), .W58(W58TO16), .W59(W59TO16), .W60(W60TO16), .W61(W61TO16), .W62(W62TO16), .W63(W63TO16)) neuron16(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out16));
neuron64in #(.W0(W0TO17), .W1(W1TO17), .W2(W2TO17), .W3(W3TO17), .W4(W4TO17), .W5(W5TO17), .W6(W6TO17), .W7(W7TO17), .W8(W8TO17), .W9(W9TO17), .W10(W10TO17), .W11(W11TO17), .W12(W12TO17), .W13(W13TO17), .W14(W14TO17), .W15(W15TO17), .W16(W16TO17), .W17(W17TO17), .W18(W18TO17), .W19(W19TO17), .W20(W20TO17), .W21(W21TO17), .W22(W22TO17), .W23(W23TO17), .W24(W24TO17), .W25(W25TO17), .W26(W26TO17), .W27(W27TO17), .W28(W28TO17), .W29(W29TO17), .W30(W30TO17), .W31(W31TO17), .W32(W32TO17), .W33(W33TO17), .W34(W34TO17), .W35(W35TO17), .W36(W36TO17), .W37(W37TO17), .W38(W38TO17), .W39(W39TO17), .W40(W40TO17), .W41(W41TO17), .W42(W42TO17), .W43(W43TO17), .W44(W44TO17), .W45(W45TO17), .W46(W46TO17), .W47(W47TO17), .W48(W48TO17), .W49(W49TO17), .W50(W50TO17), .W51(W51TO17), .W52(W52TO17), .W53(W53TO17), .W54(W54TO17), .W55(W55TO17), .W56(W56TO17), .W57(W57TO17), .W58(W58TO17), .W59(W59TO17), .W60(W60TO17), .W61(W61TO17), .W62(W62TO17), .W63(W63TO17)) neuron17(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out17));
neuron64in #(.W0(W0TO18), .W1(W1TO18), .W2(W2TO18), .W3(W3TO18), .W4(W4TO18), .W5(W5TO18), .W6(W6TO18), .W7(W7TO18), .W8(W8TO18), .W9(W9TO18), .W10(W10TO18), .W11(W11TO18), .W12(W12TO18), .W13(W13TO18), .W14(W14TO18), .W15(W15TO18), .W16(W16TO18), .W17(W17TO18), .W18(W18TO18), .W19(W19TO18), .W20(W20TO18), .W21(W21TO18), .W22(W22TO18), .W23(W23TO18), .W24(W24TO18), .W25(W25TO18), .W26(W26TO18), .W27(W27TO18), .W28(W28TO18), .W29(W29TO18), .W30(W30TO18), .W31(W31TO18), .W32(W32TO18), .W33(W33TO18), .W34(W34TO18), .W35(W35TO18), .W36(W36TO18), .W37(W37TO18), .W38(W38TO18), .W39(W39TO18), .W40(W40TO18), .W41(W41TO18), .W42(W42TO18), .W43(W43TO18), .W44(W44TO18), .W45(W45TO18), .W46(W46TO18), .W47(W47TO18), .W48(W48TO18), .W49(W49TO18), .W50(W50TO18), .W51(W51TO18), .W52(W52TO18), .W53(W53TO18), .W54(W54TO18), .W55(W55TO18), .W56(W56TO18), .W57(W57TO18), .W58(W58TO18), .W59(W59TO18), .W60(W60TO18), .W61(W61TO18), .W62(W62TO18), .W63(W63TO18)) neuron18(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out18));
neuron64in #(.W0(W0TO19), .W1(W1TO19), .W2(W2TO19), .W3(W3TO19), .W4(W4TO19), .W5(W5TO19), .W6(W6TO19), .W7(W7TO19), .W8(W8TO19), .W9(W9TO19), .W10(W10TO19), .W11(W11TO19), .W12(W12TO19), .W13(W13TO19), .W14(W14TO19), .W15(W15TO19), .W16(W16TO19), .W17(W17TO19), .W18(W18TO19), .W19(W19TO19), .W20(W20TO19), .W21(W21TO19), .W22(W22TO19), .W23(W23TO19), .W24(W24TO19), .W25(W25TO19), .W26(W26TO19), .W27(W27TO19), .W28(W28TO19), .W29(W29TO19), .W30(W30TO19), .W31(W31TO19), .W32(W32TO19), .W33(W33TO19), .W34(W34TO19), .W35(W35TO19), .W36(W36TO19), .W37(W37TO19), .W38(W38TO19), .W39(W39TO19), .W40(W40TO19), .W41(W41TO19), .W42(W42TO19), .W43(W43TO19), .W44(W44TO19), .W45(W45TO19), .W46(W46TO19), .W47(W47TO19), .W48(W48TO19), .W49(W49TO19), .W50(W50TO19), .W51(W51TO19), .W52(W52TO19), .W53(W53TO19), .W54(W54TO19), .W55(W55TO19), .W56(W56TO19), .W57(W57TO19), .W58(W58TO19), .W59(W59TO19), .W60(W60TO19), .W61(W61TO19), .W62(W62TO19), .W63(W63TO19)) neuron19(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out19));
neuron64in #(.W0(W0TO20), .W1(W1TO20), .W2(W2TO20), .W3(W3TO20), .W4(W4TO20), .W5(W5TO20), .W6(W6TO20), .W7(W7TO20), .W8(W8TO20), .W9(W9TO20), .W10(W10TO20), .W11(W11TO20), .W12(W12TO20), .W13(W13TO20), .W14(W14TO20), .W15(W15TO20), .W16(W16TO20), .W17(W17TO20), .W18(W18TO20), .W19(W19TO20), .W20(W20TO20), .W21(W21TO20), .W22(W22TO20), .W23(W23TO20), .W24(W24TO20), .W25(W25TO20), .W26(W26TO20), .W27(W27TO20), .W28(W28TO20), .W29(W29TO20), .W30(W30TO20), .W31(W31TO20), .W32(W32TO20), .W33(W33TO20), .W34(W34TO20), .W35(W35TO20), .W36(W36TO20), .W37(W37TO20), .W38(W38TO20), .W39(W39TO20), .W40(W40TO20), .W41(W41TO20), .W42(W42TO20), .W43(W43TO20), .W44(W44TO20), .W45(W45TO20), .W46(W46TO20), .W47(W47TO20), .W48(W48TO20), .W49(W49TO20), .W50(W50TO20), .W51(W51TO20), .W52(W52TO20), .W53(W53TO20), .W54(W54TO20), .W55(W55TO20), .W56(W56TO20), .W57(W57TO20), .W58(W58TO20), .W59(W59TO20), .W60(W60TO20), .W61(W61TO20), .W62(W62TO20), .W63(W63TO20)) neuron20(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out20));
neuron64in #(.W0(W0TO21), .W1(W1TO21), .W2(W2TO21), .W3(W3TO21), .W4(W4TO21), .W5(W5TO21), .W6(W6TO21), .W7(W7TO21), .W8(W8TO21), .W9(W9TO21), .W10(W10TO21), .W11(W11TO21), .W12(W12TO21), .W13(W13TO21), .W14(W14TO21), .W15(W15TO21), .W16(W16TO21), .W17(W17TO21), .W18(W18TO21), .W19(W19TO21), .W20(W20TO21), .W21(W21TO21), .W22(W22TO21), .W23(W23TO21), .W24(W24TO21), .W25(W25TO21), .W26(W26TO21), .W27(W27TO21), .W28(W28TO21), .W29(W29TO21), .W30(W30TO21), .W31(W31TO21), .W32(W32TO21), .W33(W33TO21), .W34(W34TO21), .W35(W35TO21), .W36(W36TO21), .W37(W37TO21), .W38(W38TO21), .W39(W39TO21), .W40(W40TO21), .W41(W41TO21), .W42(W42TO21), .W43(W43TO21), .W44(W44TO21), .W45(W45TO21), .W46(W46TO21), .W47(W47TO21), .W48(W48TO21), .W49(W49TO21), .W50(W50TO21), .W51(W51TO21), .W52(W52TO21), .W53(W53TO21), .W54(W54TO21), .W55(W55TO21), .W56(W56TO21), .W57(W57TO21), .W58(W58TO21), .W59(W59TO21), .W60(W60TO21), .W61(W61TO21), .W62(W62TO21), .W63(W63TO21)) neuron21(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out21));
neuron64in #(.W0(W0TO22), .W1(W1TO22), .W2(W2TO22), .W3(W3TO22), .W4(W4TO22), .W5(W5TO22), .W6(W6TO22), .W7(W7TO22), .W8(W8TO22), .W9(W9TO22), .W10(W10TO22), .W11(W11TO22), .W12(W12TO22), .W13(W13TO22), .W14(W14TO22), .W15(W15TO22), .W16(W16TO22), .W17(W17TO22), .W18(W18TO22), .W19(W19TO22), .W20(W20TO22), .W21(W21TO22), .W22(W22TO22), .W23(W23TO22), .W24(W24TO22), .W25(W25TO22), .W26(W26TO22), .W27(W27TO22), .W28(W28TO22), .W29(W29TO22), .W30(W30TO22), .W31(W31TO22), .W32(W32TO22), .W33(W33TO22), .W34(W34TO22), .W35(W35TO22), .W36(W36TO22), .W37(W37TO22), .W38(W38TO22), .W39(W39TO22), .W40(W40TO22), .W41(W41TO22), .W42(W42TO22), .W43(W43TO22), .W44(W44TO22), .W45(W45TO22), .W46(W46TO22), .W47(W47TO22), .W48(W48TO22), .W49(W49TO22), .W50(W50TO22), .W51(W51TO22), .W52(W52TO22), .W53(W53TO22), .W54(W54TO22), .W55(W55TO22), .W56(W56TO22), .W57(W57TO22), .W58(W58TO22), .W59(W59TO22), .W60(W60TO22), .W61(W61TO22), .W62(W62TO22), .W63(W63TO22)) neuron22(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out22));
neuron64in #(.W0(W0TO23), .W1(W1TO23), .W2(W2TO23), .W3(W3TO23), .W4(W4TO23), .W5(W5TO23), .W6(W6TO23), .W7(W7TO23), .W8(W8TO23), .W9(W9TO23), .W10(W10TO23), .W11(W11TO23), .W12(W12TO23), .W13(W13TO23), .W14(W14TO23), .W15(W15TO23), .W16(W16TO23), .W17(W17TO23), .W18(W18TO23), .W19(W19TO23), .W20(W20TO23), .W21(W21TO23), .W22(W22TO23), .W23(W23TO23), .W24(W24TO23), .W25(W25TO23), .W26(W26TO23), .W27(W27TO23), .W28(W28TO23), .W29(W29TO23), .W30(W30TO23), .W31(W31TO23), .W32(W32TO23), .W33(W33TO23), .W34(W34TO23), .W35(W35TO23), .W36(W36TO23), .W37(W37TO23), .W38(W38TO23), .W39(W39TO23), .W40(W40TO23), .W41(W41TO23), .W42(W42TO23), .W43(W43TO23), .W44(W44TO23), .W45(W45TO23), .W46(W46TO23), .W47(W47TO23), .W48(W48TO23), .W49(W49TO23), .W50(W50TO23), .W51(W51TO23), .W52(W52TO23), .W53(W53TO23), .W54(W54TO23), .W55(W55TO23), .W56(W56TO23), .W57(W57TO23), .W58(W58TO23), .W59(W59TO23), .W60(W60TO23), .W61(W61TO23), .W62(W62TO23), .W63(W63TO23)) neuron23(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out23));
neuron64in #(.W0(W0TO24), .W1(W1TO24), .W2(W2TO24), .W3(W3TO24), .W4(W4TO24), .W5(W5TO24), .W6(W6TO24), .W7(W7TO24), .W8(W8TO24), .W9(W9TO24), .W10(W10TO24), .W11(W11TO24), .W12(W12TO24), .W13(W13TO24), .W14(W14TO24), .W15(W15TO24), .W16(W16TO24), .W17(W17TO24), .W18(W18TO24), .W19(W19TO24), .W20(W20TO24), .W21(W21TO24), .W22(W22TO24), .W23(W23TO24), .W24(W24TO24), .W25(W25TO24), .W26(W26TO24), .W27(W27TO24), .W28(W28TO24), .W29(W29TO24), .W30(W30TO24), .W31(W31TO24), .W32(W32TO24), .W33(W33TO24), .W34(W34TO24), .W35(W35TO24), .W36(W36TO24), .W37(W37TO24), .W38(W38TO24), .W39(W39TO24), .W40(W40TO24), .W41(W41TO24), .W42(W42TO24), .W43(W43TO24), .W44(W44TO24), .W45(W45TO24), .W46(W46TO24), .W47(W47TO24), .W48(W48TO24), .W49(W49TO24), .W50(W50TO24), .W51(W51TO24), .W52(W52TO24), .W53(W53TO24), .W54(W54TO24), .W55(W55TO24), .W56(W56TO24), .W57(W57TO24), .W58(W58TO24), .W59(W59TO24), .W60(W60TO24), .W61(W61TO24), .W62(W62TO24), .W63(W63TO24)) neuron24(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out24));
neuron64in #(.W0(W0TO25), .W1(W1TO25), .W2(W2TO25), .W3(W3TO25), .W4(W4TO25), .W5(W5TO25), .W6(W6TO25), .W7(W7TO25), .W8(W8TO25), .W9(W9TO25), .W10(W10TO25), .W11(W11TO25), .W12(W12TO25), .W13(W13TO25), .W14(W14TO25), .W15(W15TO25), .W16(W16TO25), .W17(W17TO25), .W18(W18TO25), .W19(W19TO25), .W20(W20TO25), .W21(W21TO25), .W22(W22TO25), .W23(W23TO25), .W24(W24TO25), .W25(W25TO25), .W26(W26TO25), .W27(W27TO25), .W28(W28TO25), .W29(W29TO25), .W30(W30TO25), .W31(W31TO25), .W32(W32TO25), .W33(W33TO25), .W34(W34TO25), .W35(W35TO25), .W36(W36TO25), .W37(W37TO25), .W38(W38TO25), .W39(W39TO25), .W40(W40TO25), .W41(W41TO25), .W42(W42TO25), .W43(W43TO25), .W44(W44TO25), .W45(W45TO25), .W46(W46TO25), .W47(W47TO25), .W48(W48TO25), .W49(W49TO25), .W50(W50TO25), .W51(W51TO25), .W52(W52TO25), .W53(W53TO25), .W54(W54TO25), .W55(W55TO25), .W56(W56TO25), .W57(W57TO25), .W58(W58TO25), .W59(W59TO25), .W60(W60TO25), .W61(W61TO25), .W62(W62TO25), .W63(W63TO25)) neuron25(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out25));
neuron64in #(.W0(W0TO26), .W1(W1TO26), .W2(W2TO26), .W3(W3TO26), .W4(W4TO26), .W5(W5TO26), .W6(W6TO26), .W7(W7TO26), .W8(W8TO26), .W9(W9TO26), .W10(W10TO26), .W11(W11TO26), .W12(W12TO26), .W13(W13TO26), .W14(W14TO26), .W15(W15TO26), .W16(W16TO26), .W17(W17TO26), .W18(W18TO26), .W19(W19TO26), .W20(W20TO26), .W21(W21TO26), .W22(W22TO26), .W23(W23TO26), .W24(W24TO26), .W25(W25TO26), .W26(W26TO26), .W27(W27TO26), .W28(W28TO26), .W29(W29TO26), .W30(W30TO26), .W31(W31TO26), .W32(W32TO26), .W33(W33TO26), .W34(W34TO26), .W35(W35TO26), .W36(W36TO26), .W37(W37TO26), .W38(W38TO26), .W39(W39TO26), .W40(W40TO26), .W41(W41TO26), .W42(W42TO26), .W43(W43TO26), .W44(W44TO26), .W45(W45TO26), .W46(W46TO26), .W47(W47TO26), .W48(W48TO26), .W49(W49TO26), .W50(W50TO26), .W51(W51TO26), .W52(W52TO26), .W53(W53TO26), .W54(W54TO26), .W55(W55TO26), .W56(W56TO26), .W57(W57TO26), .W58(W58TO26), .W59(W59TO26), .W60(W60TO26), .W61(W61TO26), .W62(W62TO26), .W63(W63TO26)) neuron26(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out26));
neuron64in #(.W0(W0TO27), .W1(W1TO27), .W2(W2TO27), .W3(W3TO27), .W4(W4TO27), .W5(W5TO27), .W6(W6TO27), .W7(W7TO27), .W8(W8TO27), .W9(W9TO27), .W10(W10TO27), .W11(W11TO27), .W12(W12TO27), .W13(W13TO27), .W14(W14TO27), .W15(W15TO27), .W16(W16TO27), .W17(W17TO27), .W18(W18TO27), .W19(W19TO27), .W20(W20TO27), .W21(W21TO27), .W22(W22TO27), .W23(W23TO27), .W24(W24TO27), .W25(W25TO27), .W26(W26TO27), .W27(W27TO27), .W28(W28TO27), .W29(W29TO27), .W30(W30TO27), .W31(W31TO27), .W32(W32TO27), .W33(W33TO27), .W34(W34TO27), .W35(W35TO27), .W36(W36TO27), .W37(W37TO27), .W38(W38TO27), .W39(W39TO27), .W40(W40TO27), .W41(W41TO27), .W42(W42TO27), .W43(W43TO27), .W44(W44TO27), .W45(W45TO27), .W46(W46TO27), .W47(W47TO27), .W48(W48TO27), .W49(W49TO27), .W50(W50TO27), .W51(W51TO27), .W52(W52TO27), .W53(W53TO27), .W54(W54TO27), .W55(W55TO27), .W56(W56TO27), .W57(W57TO27), .W58(W58TO27), .W59(W59TO27), .W60(W60TO27), .W61(W61TO27), .W62(W62TO27), .W63(W63TO27)) neuron27(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out27));
neuron64in #(.W0(W0TO28), .W1(W1TO28), .W2(W2TO28), .W3(W3TO28), .W4(W4TO28), .W5(W5TO28), .W6(W6TO28), .W7(W7TO28), .W8(W8TO28), .W9(W9TO28), .W10(W10TO28), .W11(W11TO28), .W12(W12TO28), .W13(W13TO28), .W14(W14TO28), .W15(W15TO28), .W16(W16TO28), .W17(W17TO28), .W18(W18TO28), .W19(W19TO28), .W20(W20TO28), .W21(W21TO28), .W22(W22TO28), .W23(W23TO28), .W24(W24TO28), .W25(W25TO28), .W26(W26TO28), .W27(W27TO28), .W28(W28TO28), .W29(W29TO28), .W30(W30TO28), .W31(W31TO28), .W32(W32TO28), .W33(W33TO28), .W34(W34TO28), .W35(W35TO28), .W36(W36TO28), .W37(W37TO28), .W38(W38TO28), .W39(W39TO28), .W40(W40TO28), .W41(W41TO28), .W42(W42TO28), .W43(W43TO28), .W44(W44TO28), .W45(W45TO28), .W46(W46TO28), .W47(W47TO28), .W48(W48TO28), .W49(W49TO28), .W50(W50TO28), .W51(W51TO28), .W52(W52TO28), .W53(W53TO28), .W54(W54TO28), .W55(W55TO28), .W56(W56TO28), .W57(W57TO28), .W58(W58TO28), .W59(W59TO28), .W60(W60TO28), .W61(W61TO28), .W62(W62TO28), .W63(W63TO28)) neuron28(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out28));
neuron64in #(.W0(W0TO29), .W1(W1TO29), .W2(W2TO29), .W3(W3TO29), .W4(W4TO29), .W5(W5TO29), .W6(W6TO29), .W7(W7TO29), .W8(W8TO29), .W9(W9TO29), .W10(W10TO29), .W11(W11TO29), .W12(W12TO29), .W13(W13TO29), .W14(W14TO29), .W15(W15TO29), .W16(W16TO29), .W17(W17TO29), .W18(W18TO29), .W19(W19TO29), .W20(W20TO29), .W21(W21TO29), .W22(W22TO29), .W23(W23TO29), .W24(W24TO29), .W25(W25TO29), .W26(W26TO29), .W27(W27TO29), .W28(W28TO29), .W29(W29TO29), .W30(W30TO29), .W31(W31TO29), .W32(W32TO29), .W33(W33TO29), .W34(W34TO29), .W35(W35TO29), .W36(W36TO29), .W37(W37TO29), .W38(W38TO29), .W39(W39TO29), .W40(W40TO29), .W41(W41TO29), .W42(W42TO29), .W43(W43TO29), .W44(W44TO29), .W45(W45TO29), .W46(W46TO29), .W47(W47TO29), .W48(W48TO29), .W49(W49TO29), .W50(W50TO29), .W51(W51TO29), .W52(W52TO29), .W53(W53TO29), .W54(W54TO29), .W55(W55TO29), .W56(W56TO29), .W57(W57TO29), .W58(W58TO29), .W59(W59TO29), .W60(W60TO29), .W61(W61TO29), .W62(W62TO29), .W63(W63TO29)) neuron29(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out29));
neuron64in #(.W0(W0TO30), .W1(W1TO30), .W2(W2TO30), .W3(W3TO30), .W4(W4TO30), .W5(W5TO30), .W6(W6TO30), .W7(W7TO30), .W8(W8TO30), .W9(W9TO30), .W10(W10TO30), .W11(W11TO30), .W12(W12TO30), .W13(W13TO30), .W14(W14TO30), .W15(W15TO30), .W16(W16TO30), .W17(W17TO30), .W18(W18TO30), .W19(W19TO30), .W20(W20TO30), .W21(W21TO30), .W22(W22TO30), .W23(W23TO30), .W24(W24TO30), .W25(W25TO30), .W26(W26TO30), .W27(W27TO30), .W28(W28TO30), .W29(W29TO30), .W30(W30TO30), .W31(W31TO30), .W32(W32TO30), .W33(W33TO30), .W34(W34TO30), .W35(W35TO30), .W36(W36TO30), .W37(W37TO30), .W38(W38TO30), .W39(W39TO30), .W40(W40TO30), .W41(W41TO30), .W42(W42TO30), .W43(W43TO30), .W44(W44TO30), .W45(W45TO30), .W46(W46TO30), .W47(W47TO30), .W48(W48TO30), .W49(W49TO30), .W50(W50TO30), .W51(W51TO30), .W52(W52TO30), .W53(W53TO30), .W54(W54TO30), .W55(W55TO30), .W56(W56TO30), .W57(W57TO30), .W58(W58TO30), .W59(W59TO30), .W60(W60TO30), .W61(W61TO30), .W62(W62TO30), .W63(W63TO30)) neuron30(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out30));
neuron64in #(.W0(W0TO31), .W1(W1TO31), .W2(W2TO31), .W3(W3TO31), .W4(W4TO31), .W5(W5TO31), .W6(W6TO31), .W7(W7TO31), .W8(W8TO31), .W9(W9TO31), .W10(W10TO31), .W11(W11TO31), .W12(W12TO31), .W13(W13TO31), .W14(W14TO31), .W15(W15TO31), .W16(W16TO31), .W17(W17TO31), .W18(W18TO31), .W19(W19TO31), .W20(W20TO31), .W21(W21TO31), .W22(W22TO31), .W23(W23TO31), .W24(W24TO31), .W25(W25TO31), .W26(W26TO31), .W27(W27TO31), .W28(W28TO31), .W29(W29TO31), .W30(W30TO31), .W31(W31TO31), .W32(W32TO31), .W33(W33TO31), .W34(W34TO31), .W35(W35TO31), .W36(W36TO31), .W37(W37TO31), .W38(W38TO31), .W39(W39TO31), .W40(W40TO31), .W41(W41TO31), .W42(W42TO31), .W43(W43TO31), .W44(W44TO31), .W45(W45TO31), .W46(W46TO31), .W47(W47TO31), .W48(W48TO31), .W49(W49TO31), .W50(W50TO31), .W51(W51TO31), .W52(W52TO31), .W53(W53TO31), .W54(W54TO31), .W55(W55TO31), .W56(W56TO31), .W57(W57TO31), .W58(W58TO31), .W59(W59TO31), .W60(W60TO31), .W61(W61TO31), .W62(W62TO31), .W63(W63TO31)) neuron31(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out31));
neuron64in #(.W0(W0TO32), .W1(W1TO32), .W2(W2TO32), .W3(W3TO32), .W4(W4TO32), .W5(W5TO32), .W6(W6TO32), .W7(W7TO32), .W8(W8TO32), .W9(W9TO32), .W10(W10TO32), .W11(W11TO32), .W12(W12TO32), .W13(W13TO32), .W14(W14TO32), .W15(W15TO32), .W16(W16TO32), .W17(W17TO32), .W18(W18TO32), .W19(W19TO32), .W20(W20TO32), .W21(W21TO32), .W22(W22TO32), .W23(W23TO32), .W24(W24TO32), .W25(W25TO32), .W26(W26TO32), .W27(W27TO32), .W28(W28TO32), .W29(W29TO32), .W30(W30TO32), .W31(W31TO32), .W32(W32TO32), .W33(W33TO32), .W34(W34TO32), .W35(W35TO32), .W36(W36TO32), .W37(W37TO32), .W38(W38TO32), .W39(W39TO32), .W40(W40TO32), .W41(W41TO32), .W42(W42TO32), .W43(W43TO32), .W44(W44TO32), .W45(W45TO32), .W46(W46TO32), .W47(W47TO32), .W48(W48TO32), .W49(W49TO32), .W50(W50TO32), .W51(W51TO32), .W52(W52TO32), .W53(W53TO32), .W54(W54TO32), .W55(W55TO32), .W56(W56TO32), .W57(W57TO32), .W58(W58TO32), .W59(W59TO32), .W60(W60TO32), .W61(W61TO32), .W62(W62TO32), .W63(W63TO32)) neuron32(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out32));
neuron64in #(.W0(W0TO33), .W1(W1TO33), .W2(W2TO33), .W3(W3TO33), .W4(W4TO33), .W5(W5TO33), .W6(W6TO33), .W7(W7TO33), .W8(W8TO33), .W9(W9TO33), .W10(W10TO33), .W11(W11TO33), .W12(W12TO33), .W13(W13TO33), .W14(W14TO33), .W15(W15TO33), .W16(W16TO33), .W17(W17TO33), .W18(W18TO33), .W19(W19TO33), .W20(W20TO33), .W21(W21TO33), .W22(W22TO33), .W23(W23TO33), .W24(W24TO33), .W25(W25TO33), .W26(W26TO33), .W27(W27TO33), .W28(W28TO33), .W29(W29TO33), .W30(W30TO33), .W31(W31TO33), .W32(W32TO33), .W33(W33TO33), .W34(W34TO33), .W35(W35TO33), .W36(W36TO33), .W37(W37TO33), .W38(W38TO33), .W39(W39TO33), .W40(W40TO33), .W41(W41TO33), .W42(W42TO33), .W43(W43TO33), .W44(W44TO33), .W45(W45TO33), .W46(W46TO33), .W47(W47TO33), .W48(W48TO33), .W49(W49TO33), .W50(W50TO33), .W51(W51TO33), .W52(W52TO33), .W53(W53TO33), .W54(W54TO33), .W55(W55TO33), .W56(W56TO33), .W57(W57TO33), .W58(W58TO33), .W59(W59TO33), .W60(W60TO33), .W61(W61TO33), .W62(W62TO33), .W63(W63TO33)) neuron33(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out33));
neuron64in #(.W0(W0TO34), .W1(W1TO34), .W2(W2TO34), .W3(W3TO34), .W4(W4TO34), .W5(W5TO34), .W6(W6TO34), .W7(W7TO34), .W8(W8TO34), .W9(W9TO34), .W10(W10TO34), .W11(W11TO34), .W12(W12TO34), .W13(W13TO34), .W14(W14TO34), .W15(W15TO34), .W16(W16TO34), .W17(W17TO34), .W18(W18TO34), .W19(W19TO34), .W20(W20TO34), .W21(W21TO34), .W22(W22TO34), .W23(W23TO34), .W24(W24TO34), .W25(W25TO34), .W26(W26TO34), .W27(W27TO34), .W28(W28TO34), .W29(W29TO34), .W30(W30TO34), .W31(W31TO34), .W32(W32TO34), .W33(W33TO34), .W34(W34TO34), .W35(W35TO34), .W36(W36TO34), .W37(W37TO34), .W38(W38TO34), .W39(W39TO34), .W40(W40TO34), .W41(W41TO34), .W42(W42TO34), .W43(W43TO34), .W44(W44TO34), .W45(W45TO34), .W46(W46TO34), .W47(W47TO34), .W48(W48TO34), .W49(W49TO34), .W50(W50TO34), .W51(W51TO34), .W52(W52TO34), .W53(W53TO34), .W54(W54TO34), .W55(W55TO34), .W56(W56TO34), .W57(W57TO34), .W58(W58TO34), .W59(W59TO34), .W60(W60TO34), .W61(W61TO34), .W62(W62TO34), .W63(W63TO34)) neuron34(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out34));
neuron64in #(.W0(W0TO35), .W1(W1TO35), .W2(W2TO35), .W3(W3TO35), .W4(W4TO35), .W5(W5TO35), .W6(W6TO35), .W7(W7TO35), .W8(W8TO35), .W9(W9TO35), .W10(W10TO35), .W11(W11TO35), .W12(W12TO35), .W13(W13TO35), .W14(W14TO35), .W15(W15TO35), .W16(W16TO35), .W17(W17TO35), .W18(W18TO35), .W19(W19TO35), .W20(W20TO35), .W21(W21TO35), .W22(W22TO35), .W23(W23TO35), .W24(W24TO35), .W25(W25TO35), .W26(W26TO35), .W27(W27TO35), .W28(W28TO35), .W29(W29TO35), .W30(W30TO35), .W31(W31TO35), .W32(W32TO35), .W33(W33TO35), .W34(W34TO35), .W35(W35TO35), .W36(W36TO35), .W37(W37TO35), .W38(W38TO35), .W39(W39TO35), .W40(W40TO35), .W41(W41TO35), .W42(W42TO35), .W43(W43TO35), .W44(W44TO35), .W45(W45TO35), .W46(W46TO35), .W47(W47TO35), .W48(W48TO35), .W49(W49TO35), .W50(W50TO35), .W51(W51TO35), .W52(W52TO35), .W53(W53TO35), .W54(W54TO35), .W55(W55TO35), .W56(W56TO35), .W57(W57TO35), .W58(W58TO35), .W59(W59TO35), .W60(W60TO35), .W61(W61TO35), .W62(W62TO35), .W63(W63TO35)) neuron35(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out35));
neuron64in #(.W0(W0TO36), .W1(W1TO36), .W2(W2TO36), .W3(W3TO36), .W4(W4TO36), .W5(W5TO36), .W6(W6TO36), .W7(W7TO36), .W8(W8TO36), .W9(W9TO36), .W10(W10TO36), .W11(W11TO36), .W12(W12TO36), .W13(W13TO36), .W14(W14TO36), .W15(W15TO36), .W16(W16TO36), .W17(W17TO36), .W18(W18TO36), .W19(W19TO36), .W20(W20TO36), .W21(W21TO36), .W22(W22TO36), .W23(W23TO36), .W24(W24TO36), .W25(W25TO36), .W26(W26TO36), .W27(W27TO36), .W28(W28TO36), .W29(W29TO36), .W30(W30TO36), .W31(W31TO36), .W32(W32TO36), .W33(W33TO36), .W34(W34TO36), .W35(W35TO36), .W36(W36TO36), .W37(W37TO36), .W38(W38TO36), .W39(W39TO36), .W40(W40TO36), .W41(W41TO36), .W42(W42TO36), .W43(W43TO36), .W44(W44TO36), .W45(W45TO36), .W46(W46TO36), .W47(W47TO36), .W48(W48TO36), .W49(W49TO36), .W50(W50TO36), .W51(W51TO36), .W52(W52TO36), .W53(W53TO36), .W54(W54TO36), .W55(W55TO36), .W56(W56TO36), .W57(W57TO36), .W58(W58TO36), .W59(W59TO36), .W60(W60TO36), .W61(W61TO36), .W62(W62TO36), .W63(W63TO36)) neuron36(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out36));
neuron64in #(.W0(W0TO37), .W1(W1TO37), .W2(W2TO37), .W3(W3TO37), .W4(W4TO37), .W5(W5TO37), .W6(W6TO37), .W7(W7TO37), .W8(W8TO37), .W9(W9TO37), .W10(W10TO37), .W11(W11TO37), .W12(W12TO37), .W13(W13TO37), .W14(W14TO37), .W15(W15TO37), .W16(W16TO37), .W17(W17TO37), .W18(W18TO37), .W19(W19TO37), .W20(W20TO37), .W21(W21TO37), .W22(W22TO37), .W23(W23TO37), .W24(W24TO37), .W25(W25TO37), .W26(W26TO37), .W27(W27TO37), .W28(W28TO37), .W29(W29TO37), .W30(W30TO37), .W31(W31TO37), .W32(W32TO37), .W33(W33TO37), .W34(W34TO37), .W35(W35TO37), .W36(W36TO37), .W37(W37TO37), .W38(W38TO37), .W39(W39TO37), .W40(W40TO37), .W41(W41TO37), .W42(W42TO37), .W43(W43TO37), .W44(W44TO37), .W45(W45TO37), .W46(W46TO37), .W47(W47TO37), .W48(W48TO37), .W49(W49TO37), .W50(W50TO37), .W51(W51TO37), .W52(W52TO37), .W53(W53TO37), .W54(W54TO37), .W55(W55TO37), .W56(W56TO37), .W57(W57TO37), .W58(W58TO37), .W59(W59TO37), .W60(W60TO37), .W61(W61TO37), .W62(W62TO37), .W63(W63TO37)) neuron37(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out37));
neuron64in #(.W0(W0TO38), .W1(W1TO38), .W2(W2TO38), .W3(W3TO38), .W4(W4TO38), .W5(W5TO38), .W6(W6TO38), .W7(W7TO38), .W8(W8TO38), .W9(W9TO38), .W10(W10TO38), .W11(W11TO38), .W12(W12TO38), .W13(W13TO38), .W14(W14TO38), .W15(W15TO38), .W16(W16TO38), .W17(W17TO38), .W18(W18TO38), .W19(W19TO38), .W20(W20TO38), .W21(W21TO38), .W22(W22TO38), .W23(W23TO38), .W24(W24TO38), .W25(W25TO38), .W26(W26TO38), .W27(W27TO38), .W28(W28TO38), .W29(W29TO38), .W30(W30TO38), .W31(W31TO38), .W32(W32TO38), .W33(W33TO38), .W34(W34TO38), .W35(W35TO38), .W36(W36TO38), .W37(W37TO38), .W38(W38TO38), .W39(W39TO38), .W40(W40TO38), .W41(W41TO38), .W42(W42TO38), .W43(W43TO38), .W44(W44TO38), .W45(W45TO38), .W46(W46TO38), .W47(W47TO38), .W48(W48TO38), .W49(W49TO38), .W50(W50TO38), .W51(W51TO38), .W52(W52TO38), .W53(W53TO38), .W54(W54TO38), .W55(W55TO38), .W56(W56TO38), .W57(W57TO38), .W58(W58TO38), .W59(W59TO38), .W60(W60TO38), .W61(W61TO38), .W62(W62TO38), .W63(W63TO38)) neuron38(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out38));
neuron64in #(.W0(W0TO39), .W1(W1TO39), .W2(W2TO39), .W3(W3TO39), .W4(W4TO39), .W5(W5TO39), .W6(W6TO39), .W7(W7TO39), .W8(W8TO39), .W9(W9TO39), .W10(W10TO39), .W11(W11TO39), .W12(W12TO39), .W13(W13TO39), .W14(W14TO39), .W15(W15TO39), .W16(W16TO39), .W17(W17TO39), .W18(W18TO39), .W19(W19TO39), .W20(W20TO39), .W21(W21TO39), .W22(W22TO39), .W23(W23TO39), .W24(W24TO39), .W25(W25TO39), .W26(W26TO39), .W27(W27TO39), .W28(W28TO39), .W29(W29TO39), .W30(W30TO39), .W31(W31TO39), .W32(W32TO39), .W33(W33TO39), .W34(W34TO39), .W35(W35TO39), .W36(W36TO39), .W37(W37TO39), .W38(W38TO39), .W39(W39TO39), .W40(W40TO39), .W41(W41TO39), .W42(W42TO39), .W43(W43TO39), .W44(W44TO39), .W45(W45TO39), .W46(W46TO39), .W47(W47TO39), .W48(W48TO39), .W49(W49TO39), .W50(W50TO39), .W51(W51TO39), .W52(W52TO39), .W53(W53TO39), .W54(W54TO39), .W55(W55TO39), .W56(W56TO39), .W57(W57TO39), .W58(W58TO39), .W59(W59TO39), .W60(W60TO39), .W61(W61TO39), .W62(W62TO39), .W63(W63TO39)) neuron39(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out39));
neuron64in #(.W0(W0TO40), .W1(W1TO40), .W2(W2TO40), .W3(W3TO40), .W4(W4TO40), .W5(W5TO40), .W6(W6TO40), .W7(W7TO40), .W8(W8TO40), .W9(W9TO40), .W10(W10TO40), .W11(W11TO40), .W12(W12TO40), .W13(W13TO40), .W14(W14TO40), .W15(W15TO40), .W16(W16TO40), .W17(W17TO40), .W18(W18TO40), .W19(W19TO40), .W20(W20TO40), .W21(W21TO40), .W22(W22TO40), .W23(W23TO40), .W24(W24TO40), .W25(W25TO40), .W26(W26TO40), .W27(W27TO40), .W28(W28TO40), .W29(W29TO40), .W30(W30TO40), .W31(W31TO40), .W32(W32TO40), .W33(W33TO40), .W34(W34TO40), .W35(W35TO40), .W36(W36TO40), .W37(W37TO40), .W38(W38TO40), .W39(W39TO40), .W40(W40TO40), .W41(W41TO40), .W42(W42TO40), .W43(W43TO40), .W44(W44TO40), .W45(W45TO40), .W46(W46TO40), .W47(W47TO40), .W48(W48TO40), .W49(W49TO40), .W50(W50TO40), .W51(W51TO40), .W52(W52TO40), .W53(W53TO40), .W54(W54TO40), .W55(W55TO40), .W56(W56TO40), .W57(W57TO40), .W58(W58TO40), .W59(W59TO40), .W60(W60TO40), .W61(W61TO40), .W62(W62TO40), .W63(W63TO40)) neuron40(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out40));
neuron64in #(.W0(W0TO41), .W1(W1TO41), .W2(W2TO41), .W3(W3TO41), .W4(W4TO41), .W5(W5TO41), .W6(W6TO41), .W7(W7TO41), .W8(W8TO41), .W9(W9TO41), .W10(W10TO41), .W11(W11TO41), .W12(W12TO41), .W13(W13TO41), .W14(W14TO41), .W15(W15TO41), .W16(W16TO41), .W17(W17TO41), .W18(W18TO41), .W19(W19TO41), .W20(W20TO41), .W21(W21TO41), .W22(W22TO41), .W23(W23TO41), .W24(W24TO41), .W25(W25TO41), .W26(W26TO41), .W27(W27TO41), .W28(W28TO41), .W29(W29TO41), .W30(W30TO41), .W31(W31TO41), .W32(W32TO41), .W33(W33TO41), .W34(W34TO41), .W35(W35TO41), .W36(W36TO41), .W37(W37TO41), .W38(W38TO41), .W39(W39TO41), .W40(W40TO41), .W41(W41TO41), .W42(W42TO41), .W43(W43TO41), .W44(W44TO41), .W45(W45TO41), .W46(W46TO41), .W47(W47TO41), .W48(W48TO41), .W49(W49TO41), .W50(W50TO41), .W51(W51TO41), .W52(W52TO41), .W53(W53TO41), .W54(W54TO41), .W55(W55TO41), .W56(W56TO41), .W57(W57TO41), .W58(W58TO41), .W59(W59TO41), .W60(W60TO41), .W61(W61TO41), .W62(W62TO41), .W63(W63TO41)) neuron41(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out41));
neuron64in #(.W0(W0TO42), .W1(W1TO42), .W2(W2TO42), .W3(W3TO42), .W4(W4TO42), .W5(W5TO42), .W6(W6TO42), .W7(W7TO42), .W8(W8TO42), .W9(W9TO42), .W10(W10TO42), .W11(W11TO42), .W12(W12TO42), .W13(W13TO42), .W14(W14TO42), .W15(W15TO42), .W16(W16TO42), .W17(W17TO42), .W18(W18TO42), .W19(W19TO42), .W20(W20TO42), .W21(W21TO42), .W22(W22TO42), .W23(W23TO42), .W24(W24TO42), .W25(W25TO42), .W26(W26TO42), .W27(W27TO42), .W28(W28TO42), .W29(W29TO42), .W30(W30TO42), .W31(W31TO42), .W32(W32TO42), .W33(W33TO42), .W34(W34TO42), .W35(W35TO42), .W36(W36TO42), .W37(W37TO42), .W38(W38TO42), .W39(W39TO42), .W40(W40TO42), .W41(W41TO42), .W42(W42TO42), .W43(W43TO42), .W44(W44TO42), .W45(W45TO42), .W46(W46TO42), .W47(W47TO42), .W48(W48TO42), .W49(W49TO42), .W50(W50TO42), .W51(W51TO42), .W52(W52TO42), .W53(W53TO42), .W54(W54TO42), .W55(W55TO42), .W56(W56TO42), .W57(W57TO42), .W58(W58TO42), .W59(W59TO42), .W60(W60TO42), .W61(W61TO42), .W62(W62TO42), .W63(W63TO42)) neuron42(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out42));
neuron64in #(.W0(W0TO43), .W1(W1TO43), .W2(W2TO43), .W3(W3TO43), .W4(W4TO43), .W5(W5TO43), .W6(W6TO43), .W7(W7TO43), .W8(W8TO43), .W9(W9TO43), .W10(W10TO43), .W11(W11TO43), .W12(W12TO43), .W13(W13TO43), .W14(W14TO43), .W15(W15TO43), .W16(W16TO43), .W17(W17TO43), .W18(W18TO43), .W19(W19TO43), .W20(W20TO43), .W21(W21TO43), .W22(W22TO43), .W23(W23TO43), .W24(W24TO43), .W25(W25TO43), .W26(W26TO43), .W27(W27TO43), .W28(W28TO43), .W29(W29TO43), .W30(W30TO43), .W31(W31TO43), .W32(W32TO43), .W33(W33TO43), .W34(W34TO43), .W35(W35TO43), .W36(W36TO43), .W37(W37TO43), .W38(W38TO43), .W39(W39TO43), .W40(W40TO43), .W41(W41TO43), .W42(W42TO43), .W43(W43TO43), .W44(W44TO43), .W45(W45TO43), .W46(W46TO43), .W47(W47TO43), .W48(W48TO43), .W49(W49TO43), .W50(W50TO43), .W51(W51TO43), .W52(W52TO43), .W53(W53TO43), .W54(W54TO43), .W55(W55TO43), .W56(W56TO43), .W57(W57TO43), .W58(W58TO43), .W59(W59TO43), .W60(W60TO43), .W61(W61TO43), .W62(W62TO43), .W63(W63TO43)) neuron43(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out43));
neuron64in #(.W0(W0TO44), .W1(W1TO44), .W2(W2TO44), .W3(W3TO44), .W4(W4TO44), .W5(W5TO44), .W6(W6TO44), .W7(W7TO44), .W8(W8TO44), .W9(W9TO44), .W10(W10TO44), .W11(W11TO44), .W12(W12TO44), .W13(W13TO44), .W14(W14TO44), .W15(W15TO44), .W16(W16TO44), .W17(W17TO44), .W18(W18TO44), .W19(W19TO44), .W20(W20TO44), .W21(W21TO44), .W22(W22TO44), .W23(W23TO44), .W24(W24TO44), .W25(W25TO44), .W26(W26TO44), .W27(W27TO44), .W28(W28TO44), .W29(W29TO44), .W30(W30TO44), .W31(W31TO44), .W32(W32TO44), .W33(W33TO44), .W34(W34TO44), .W35(W35TO44), .W36(W36TO44), .W37(W37TO44), .W38(W38TO44), .W39(W39TO44), .W40(W40TO44), .W41(W41TO44), .W42(W42TO44), .W43(W43TO44), .W44(W44TO44), .W45(W45TO44), .W46(W46TO44), .W47(W47TO44), .W48(W48TO44), .W49(W49TO44), .W50(W50TO44), .W51(W51TO44), .W52(W52TO44), .W53(W53TO44), .W54(W54TO44), .W55(W55TO44), .W56(W56TO44), .W57(W57TO44), .W58(W58TO44), .W59(W59TO44), .W60(W60TO44), .W61(W61TO44), .W62(W62TO44), .W63(W63TO44)) neuron44(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out44));
neuron64in #(.W0(W0TO45), .W1(W1TO45), .W2(W2TO45), .W3(W3TO45), .W4(W4TO45), .W5(W5TO45), .W6(W6TO45), .W7(W7TO45), .W8(W8TO45), .W9(W9TO45), .W10(W10TO45), .W11(W11TO45), .W12(W12TO45), .W13(W13TO45), .W14(W14TO45), .W15(W15TO45), .W16(W16TO45), .W17(W17TO45), .W18(W18TO45), .W19(W19TO45), .W20(W20TO45), .W21(W21TO45), .W22(W22TO45), .W23(W23TO45), .W24(W24TO45), .W25(W25TO45), .W26(W26TO45), .W27(W27TO45), .W28(W28TO45), .W29(W29TO45), .W30(W30TO45), .W31(W31TO45), .W32(W32TO45), .W33(W33TO45), .W34(W34TO45), .W35(W35TO45), .W36(W36TO45), .W37(W37TO45), .W38(W38TO45), .W39(W39TO45), .W40(W40TO45), .W41(W41TO45), .W42(W42TO45), .W43(W43TO45), .W44(W44TO45), .W45(W45TO45), .W46(W46TO45), .W47(W47TO45), .W48(W48TO45), .W49(W49TO45), .W50(W50TO45), .W51(W51TO45), .W52(W52TO45), .W53(W53TO45), .W54(W54TO45), .W55(W55TO45), .W56(W56TO45), .W57(W57TO45), .W58(W58TO45), .W59(W59TO45), .W60(W60TO45), .W61(W61TO45), .W62(W62TO45), .W63(W63TO45)) neuron45(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out45));
neuron64in #(.W0(W0TO46), .W1(W1TO46), .W2(W2TO46), .W3(W3TO46), .W4(W4TO46), .W5(W5TO46), .W6(W6TO46), .W7(W7TO46), .W8(W8TO46), .W9(W9TO46), .W10(W10TO46), .W11(W11TO46), .W12(W12TO46), .W13(W13TO46), .W14(W14TO46), .W15(W15TO46), .W16(W16TO46), .W17(W17TO46), .W18(W18TO46), .W19(W19TO46), .W20(W20TO46), .W21(W21TO46), .W22(W22TO46), .W23(W23TO46), .W24(W24TO46), .W25(W25TO46), .W26(W26TO46), .W27(W27TO46), .W28(W28TO46), .W29(W29TO46), .W30(W30TO46), .W31(W31TO46), .W32(W32TO46), .W33(W33TO46), .W34(W34TO46), .W35(W35TO46), .W36(W36TO46), .W37(W37TO46), .W38(W38TO46), .W39(W39TO46), .W40(W40TO46), .W41(W41TO46), .W42(W42TO46), .W43(W43TO46), .W44(W44TO46), .W45(W45TO46), .W46(W46TO46), .W47(W47TO46), .W48(W48TO46), .W49(W49TO46), .W50(W50TO46), .W51(W51TO46), .W52(W52TO46), .W53(W53TO46), .W54(W54TO46), .W55(W55TO46), .W56(W56TO46), .W57(W57TO46), .W58(W58TO46), .W59(W59TO46), .W60(W60TO46), .W61(W61TO46), .W62(W62TO46), .W63(W63TO46)) neuron46(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out46));
neuron64in #(.W0(W0TO47), .W1(W1TO47), .W2(W2TO47), .W3(W3TO47), .W4(W4TO47), .W5(W5TO47), .W6(W6TO47), .W7(W7TO47), .W8(W8TO47), .W9(W9TO47), .W10(W10TO47), .W11(W11TO47), .W12(W12TO47), .W13(W13TO47), .W14(W14TO47), .W15(W15TO47), .W16(W16TO47), .W17(W17TO47), .W18(W18TO47), .W19(W19TO47), .W20(W20TO47), .W21(W21TO47), .W22(W22TO47), .W23(W23TO47), .W24(W24TO47), .W25(W25TO47), .W26(W26TO47), .W27(W27TO47), .W28(W28TO47), .W29(W29TO47), .W30(W30TO47), .W31(W31TO47), .W32(W32TO47), .W33(W33TO47), .W34(W34TO47), .W35(W35TO47), .W36(W36TO47), .W37(W37TO47), .W38(W38TO47), .W39(W39TO47), .W40(W40TO47), .W41(W41TO47), .W42(W42TO47), .W43(W43TO47), .W44(W44TO47), .W45(W45TO47), .W46(W46TO47), .W47(W47TO47), .W48(W48TO47), .W49(W49TO47), .W50(W50TO47), .W51(W51TO47), .W52(W52TO47), .W53(W53TO47), .W54(W54TO47), .W55(W55TO47), .W56(W56TO47), .W57(W57TO47), .W58(W58TO47), .W59(W59TO47), .W60(W60TO47), .W61(W61TO47), .W62(W62TO47), .W63(W63TO47)) neuron47(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out47));
neuron64in #(.W0(W0TO48), .W1(W1TO48), .W2(W2TO48), .W3(W3TO48), .W4(W4TO48), .W5(W5TO48), .W6(W6TO48), .W7(W7TO48), .W8(W8TO48), .W9(W9TO48), .W10(W10TO48), .W11(W11TO48), .W12(W12TO48), .W13(W13TO48), .W14(W14TO48), .W15(W15TO48), .W16(W16TO48), .W17(W17TO48), .W18(W18TO48), .W19(W19TO48), .W20(W20TO48), .W21(W21TO48), .W22(W22TO48), .W23(W23TO48), .W24(W24TO48), .W25(W25TO48), .W26(W26TO48), .W27(W27TO48), .W28(W28TO48), .W29(W29TO48), .W30(W30TO48), .W31(W31TO48), .W32(W32TO48), .W33(W33TO48), .W34(W34TO48), .W35(W35TO48), .W36(W36TO48), .W37(W37TO48), .W38(W38TO48), .W39(W39TO48), .W40(W40TO48), .W41(W41TO48), .W42(W42TO48), .W43(W43TO48), .W44(W44TO48), .W45(W45TO48), .W46(W46TO48), .W47(W47TO48), .W48(W48TO48), .W49(W49TO48), .W50(W50TO48), .W51(W51TO48), .W52(W52TO48), .W53(W53TO48), .W54(W54TO48), .W55(W55TO48), .W56(W56TO48), .W57(W57TO48), .W58(W58TO48), .W59(W59TO48), .W60(W60TO48), .W61(W61TO48), .W62(W62TO48), .W63(W63TO48)) neuron48(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out48));
neuron64in #(.W0(W0TO49), .W1(W1TO49), .W2(W2TO49), .W3(W3TO49), .W4(W4TO49), .W5(W5TO49), .W6(W6TO49), .W7(W7TO49), .W8(W8TO49), .W9(W9TO49), .W10(W10TO49), .W11(W11TO49), .W12(W12TO49), .W13(W13TO49), .W14(W14TO49), .W15(W15TO49), .W16(W16TO49), .W17(W17TO49), .W18(W18TO49), .W19(W19TO49), .W20(W20TO49), .W21(W21TO49), .W22(W22TO49), .W23(W23TO49), .W24(W24TO49), .W25(W25TO49), .W26(W26TO49), .W27(W27TO49), .W28(W28TO49), .W29(W29TO49), .W30(W30TO49), .W31(W31TO49), .W32(W32TO49), .W33(W33TO49), .W34(W34TO49), .W35(W35TO49), .W36(W36TO49), .W37(W37TO49), .W38(W38TO49), .W39(W39TO49), .W40(W40TO49), .W41(W41TO49), .W42(W42TO49), .W43(W43TO49), .W44(W44TO49), .W45(W45TO49), .W46(W46TO49), .W47(W47TO49), .W48(W48TO49), .W49(W49TO49), .W50(W50TO49), .W51(W51TO49), .W52(W52TO49), .W53(W53TO49), .W54(W54TO49), .W55(W55TO49), .W56(W56TO49), .W57(W57TO49), .W58(W58TO49), .W59(W59TO49), .W60(W60TO49), .W61(W61TO49), .W62(W62TO49), .W63(W63TO49)) neuron49(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out49));
neuron64in #(.W0(W0TO50), .W1(W1TO50), .W2(W2TO50), .W3(W3TO50), .W4(W4TO50), .W5(W5TO50), .W6(W6TO50), .W7(W7TO50), .W8(W8TO50), .W9(W9TO50), .W10(W10TO50), .W11(W11TO50), .W12(W12TO50), .W13(W13TO50), .W14(W14TO50), .W15(W15TO50), .W16(W16TO50), .W17(W17TO50), .W18(W18TO50), .W19(W19TO50), .W20(W20TO50), .W21(W21TO50), .W22(W22TO50), .W23(W23TO50), .W24(W24TO50), .W25(W25TO50), .W26(W26TO50), .W27(W27TO50), .W28(W28TO50), .W29(W29TO50), .W30(W30TO50), .W31(W31TO50), .W32(W32TO50), .W33(W33TO50), .W34(W34TO50), .W35(W35TO50), .W36(W36TO50), .W37(W37TO50), .W38(W38TO50), .W39(W39TO50), .W40(W40TO50), .W41(W41TO50), .W42(W42TO50), .W43(W43TO50), .W44(W44TO50), .W45(W45TO50), .W46(W46TO50), .W47(W47TO50), .W48(W48TO50), .W49(W49TO50), .W50(W50TO50), .W51(W51TO50), .W52(W52TO50), .W53(W53TO50), .W54(W54TO50), .W55(W55TO50), .W56(W56TO50), .W57(W57TO50), .W58(W58TO50), .W59(W59TO50), .W60(W60TO50), .W61(W61TO50), .W62(W62TO50), .W63(W63TO50)) neuron50(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out50));
neuron64in #(.W0(W0TO51), .W1(W1TO51), .W2(W2TO51), .W3(W3TO51), .W4(W4TO51), .W5(W5TO51), .W6(W6TO51), .W7(W7TO51), .W8(W8TO51), .W9(W9TO51), .W10(W10TO51), .W11(W11TO51), .W12(W12TO51), .W13(W13TO51), .W14(W14TO51), .W15(W15TO51), .W16(W16TO51), .W17(W17TO51), .W18(W18TO51), .W19(W19TO51), .W20(W20TO51), .W21(W21TO51), .W22(W22TO51), .W23(W23TO51), .W24(W24TO51), .W25(W25TO51), .W26(W26TO51), .W27(W27TO51), .W28(W28TO51), .W29(W29TO51), .W30(W30TO51), .W31(W31TO51), .W32(W32TO51), .W33(W33TO51), .W34(W34TO51), .W35(W35TO51), .W36(W36TO51), .W37(W37TO51), .W38(W38TO51), .W39(W39TO51), .W40(W40TO51), .W41(W41TO51), .W42(W42TO51), .W43(W43TO51), .W44(W44TO51), .W45(W45TO51), .W46(W46TO51), .W47(W47TO51), .W48(W48TO51), .W49(W49TO51), .W50(W50TO51), .W51(W51TO51), .W52(W52TO51), .W53(W53TO51), .W54(W54TO51), .W55(W55TO51), .W56(W56TO51), .W57(W57TO51), .W58(W58TO51), .W59(W59TO51), .W60(W60TO51), .W61(W61TO51), .W62(W62TO51), .W63(W63TO51)) neuron51(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out51));
neuron64in #(.W0(W0TO52), .W1(W1TO52), .W2(W2TO52), .W3(W3TO52), .W4(W4TO52), .W5(W5TO52), .W6(W6TO52), .W7(W7TO52), .W8(W8TO52), .W9(W9TO52), .W10(W10TO52), .W11(W11TO52), .W12(W12TO52), .W13(W13TO52), .W14(W14TO52), .W15(W15TO52), .W16(W16TO52), .W17(W17TO52), .W18(W18TO52), .W19(W19TO52), .W20(W20TO52), .W21(W21TO52), .W22(W22TO52), .W23(W23TO52), .W24(W24TO52), .W25(W25TO52), .W26(W26TO52), .W27(W27TO52), .W28(W28TO52), .W29(W29TO52), .W30(W30TO52), .W31(W31TO52), .W32(W32TO52), .W33(W33TO52), .W34(W34TO52), .W35(W35TO52), .W36(W36TO52), .W37(W37TO52), .W38(W38TO52), .W39(W39TO52), .W40(W40TO52), .W41(W41TO52), .W42(W42TO52), .W43(W43TO52), .W44(W44TO52), .W45(W45TO52), .W46(W46TO52), .W47(W47TO52), .W48(W48TO52), .W49(W49TO52), .W50(W50TO52), .W51(W51TO52), .W52(W52TO52), .W53(W53TO52), .W54(W54TO52), .W55(W55TO52), .W56(W56TO52), .W57(W57TO52), .W58(W58TO52), .W59(W59TO52), .W60(W60TO52), .W61(W61TO52), .W62(W62TO52), .W63(W63TO52)) neuron52(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out52));
neuron64in #(.W0(W0TO53), .W1(W1TO53), .W2(W2TO53), .W3(W3TO53), .W4(W4TO53), .W5(W5TO53), .W6(W6TO53), .W7(W7TO53), .W8(W8TO53), .W9(W9TO53), .W10(W10TO53), .W11(W11TO53), .W12(W12TO53), .W13(W13TO53), .W14(W14TO53), .W15(W15TO53), .W16(W16TO53), .W17(W17TO53), .W18(W18TO53), .W19(W19TO53), .W20(W20TO53), .W21(W21TO53), .W22(W22TO53), .W23(W23TO53), .W24(W24TO53), .W25(W25TO53), .W26(W26TO53), .W27(W27TO53), .W28(W28TO53), .W29(W29TO53), .W30(W30TO53), .W31(W31TO53), .W32(W32TO53), .W33(W33TO53), .W34(W34TO53), .W35(W35TO53), .W36(W36TO53), .W37(W37TO53), .W38(W38TO53), .W39(W39TO53), .W40(W40TO53), .W41(W41TO53), .W42(W42TO53), .W43(W43TO53), .W44(W44TO53), .W45(W45TO53), .W46(W46TO53), .W47(W47TO53), .W48(W48TO53), .W49(W49TO53), .W50(W50TO53), .W51(W51TO53), .W52(W52TO53), .W53(W53TO53), .W54(W54TO53), .W55(W55TO53), .W56(W56TO53), .W57(W57TO53), .W58(W58TO53), .W59(W59TO53), .W60(W60TO53), .W61(W61TO53), .W62(W62TO53), .W63(W63TO53)) neuron53(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out53));
neuron64in #(.W0(W0TO54), .W1(W1TO54), .W2(W2TO54), .W3(W3TO54), .W4(W4TO54), .W5(W5TO54), .W6(W6TO54), .W7(W7TO54), .W8(W8TO54), .W9(W9TO54), .W10(W10TO54), .W11(W11TO54), .W12(W12TO54), .W13(W13TO54), .W14(W14TO54), .W15(W15TO54), .W16(W16TO54), .W17(W17TO54), .W18(W18TO54), .W19(W19TO54), .W20(W20TO54), .W21(W21TO54), .W22(W22TO54), .W23(W23TO54), .W24(W24TO54), .W25(W25TO54), .W26(W26TO54), .W27(W27TO54), .W28(W28TO54), .W29(W29TO54), .W30(W30TO54), .W31(W31TO54), .W32(W32TO54), .W33(W33TO54), .W34(W34TO54), .W35(W35TO54), .W36(W36TO54), .W37(W37TO54), .W38(W38TO54), .W39(W39TO54), .W40(W40TO54), .W41(W41TO54), .W42(W42TO54), .W43(W43TO54), .W44(W44TO54), .W45(W45TO54), .W46(W46TO54), .W47(W47TO54), .W48(W48TO54), .W49(W49TO54), .W50(W50TO54), .W51(W51TO54), .W52(W52TO54), .W53(W53TO54), .W54(W54TO54), .W55(W55TO54), .W56(W56TO54), .W57(W57TO54), .W58(W58TO54), .W59(W59TO54), .W60(W60TO54), .W61(W61TO54), .W62(W62TO54), .W63(W63TO54)) neuron54(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out54));
neuron64in #(.W0(W0TO55), .W1(W1TO55), .W2(W2TO55), .W3(W3TO55), .W4(W4TO55), .W5(W5TO55), .W6(W6TO55), .W7(W7TO55), .W8(W8TO55), .W9(W9TO55), .W10(W10TO55), .W11(W11TO55), .W12(W12TO55), .W13(W13TO55), .W14(W14TO55), .W15(W15TO55), .W16(W16TO55), .W17(W17TO55), .W18(W18TO55), .W19(W19TO55), .W20(W20TO55), .W21(W21TO55), .W22(W22TO55), .W23(W23TO55), .W24(W24TO55), .W25(W25TO55), .W26(W26TO55), .W27(W27TO55), .W28(W28TO55), .W29(W29TO55), .W30(W30TO55), .W31(W31TO55), .W32(W32TO55), .W33(W33TO55), .W34(W34TO55), .W35(W35TO55), .W36(W36TO55), .W37(W37TO55), .W38(W38TO55), .W39(W39TO55), .W40(W40TO55), .W41(W41TO55), .W42(W42TO55), .W43(W43TO55), .W44(W44TO55), .W45(W45TO55), .W46(W46TO55), .W47(W47TO55), .W48(W48TO55), .W49(W49TO55), .W50(W50TO55), .W51(W51TO55), .W52(W52TO55), .W53(W53TO55), .W54(W54TO55), .W55(W55TO55), .W56(W56TO55), .W57(W57TO55), .W58(W58TO55), .W59(W59TO55), .W60(W60TO55), .W61(W61TO55), .W62(W62TO55), .W63(W63TO55)) neuron55(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out55));
neuron64in #(.W0(W0TO56), .W1(W1TO56), .W2(W2TO56), .W3(W3TO56), .W4(W4TO56), .W5(W5TO56), .W6(W6TO56), .W7(W7TO56), .W8(W8TO56), .W9(W9TO56), .W10(W10TO56), .W11(W11TO56), .W12(W12TO56), .W13(W13TO56), .W14(W14TO56), .W15(W15TO56), .W16(W16TO56), .W17(W17TO56), .W18(W18TO56), .W19(W19TO56), .W20(W20TO56), .W21(W21TO56), .W22(W22TO56), .W23(W23TO56), .W24(W24TO56), .W25(W25TO56), .W26(W26TO56), .W27(W27TO56), .W28(W28TO56), .W29(W29TO56), .W30(W30TO56), .W31(W31TO56), .W32(W32TO56), .W33(W33TO56), .W34(W34TO56), .W35(W35TO56), .W36(W36TO56), .W37(W37TO56), .W38(W38TO56), .W39(W39TO56), .W40(W40TO56), .W41(W41TO56), .W42(W42TO56), .W43(W43TO56), .W44(W44TO56), .W45(W45TO56), .W46(W46TO56), .W47(W47TO56), .W48(W48TO56), .W49(W49TO56), .W50(W50TO56), .W51(W51TO56), .W52(W52TO56), .W53(W53TO56), .W54(W54TO56), .W55(W55TO56), .W56(W56TO56), .W57(W57TO56), .W58(W58TO56), .W59(W59TO56), .W60(W60TO56), .W61(W61TO56), .W62(W62TO56), .W63(W63TO56)) neuron56(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out56));
neuron64in #(.W0(W0TO57), .W1(W1TO57), .W2(W2TO57), .W3(W3TO57), .W4(W4TO57), .W5(W5TO57), .W6(W6TO57), .W7(W7TO57), .W8(W8TO57), .W9(W9TO57), .W10(W10TO57), .W11(W11TO57), .W12(W12TO57), .W13(W13TO57), .W14(W14TO57), .W15(W15TO57), .W16(W16TO57), .W17(W17TO57), .W18(W18TO57), .W19(W19TO57), .W20(W20TO57), .W21(W21TO57), .W22(W22TO57), .W23(W23TO57), .W24(W24TO57), .W25(W25TO57), .W26(W26TO57), .W27(W27TO57), .W28(W28TO57), .W29(W29TO57), .W30(W30TO57), .W31(W31TO57), .W32(W32TO57), .W33(W33TO57), .W34(W34TO57), .W35(W35TO57), .W36(W36TO57), .W37(W37TO57), .W38(W38TO57), .W39(W39TO57), .W40(W40TO57), .W41(W41TO57), .W42(W42TO57), .W43(W43TO57), .W44(W44TO57), .W45(W45TO57), .W46(W46TO57), .W47(W47TO57), .W48(W48TO57), .W49(W49TO57), .W50(W50TO57), .W51(W51TO57), .W52(W52TO57), .W53(W53TO57), .W54(W54TO57), .W55(W55TO57), .W56(W56TO57), .W57(W57TO57), .W58(W58TO57), .W59(W59TO57), .W60(W60TO57), .W61(W61TO57), .W62(W62TO57), .W63(W63TO57)) neuron57(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out57));
neuron64in #(.W0(W0TO58), .W1(W1TO58), .W2(W2TO58), .W3(W3TO58), .W4(W4TO58), .W5(W5TO58), .W6(W6TO58), .W7(W7TO58), .W8(W8TO58), .W9(W9TO58), .W10(W10TO58), .W11(W11TO58), .W12(W12TO58), .W13(W13TO58), .W14(W14TO58), .W15(W15TO58), .W16(W16TO58), .W17(W17TO58), .W18(W18TO58), .W19(W19TO58), .W20(W20TO58), .W21(W21TO58), .W22(W22TO58), .W23(W23TO58), .W24(W24TO58), .W25(W25TO58), .W26(W26TO58), .W27(W27TO58), .W28(W28TO58), .W29(W29TO58), .W30(W30TO58), .W31(W31TO58), .W32(W32TO58), .W33(W33TO58), .W34(W34TO58), .W35(W35TO58), .W36(W36TO58), .W37(W37TO58), .W38(W38TO58), .W39(W39TO58), .W40(W40TO58), .W41(W41TO58), .W42(W42TO58), .W43(W43TO58), .W44(W44TO58), .W45(W45TO58), .W46(W46TO58), .W47(W47TO58), .W48(W48TO58), .W49(W49TO58), .W50(W50TO58), .W51(W51TO58), .W52(W52TO58), .W53(W53TO58), .W54(W54TO58), .W55(W55TO58), .W56(W56TO58), .W57(W57TO58), .W58(W58TO58), .W59(W59TO58), .W60(W60TO58), .W61(W61TO58), .W62(W62TO58), .W63(W63TO58)) neuron58(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out58));
neuron64in #(.W0(W0TO59), .W1(W1TO59), .W2(W2TO59), .W3(W3TO59), .W4(W4TO59), .W5(W5TO59), .W6(W6TO59), .W7(W7TO59), .W8(W8TO59), .W9(W9TO59), .W10(W10TO59), .W11(W11TO59), .W12(W12TO59), .W13(W13TO59), .W14(W14TO59), .W15(W15TO59), .W16(W16TO59), .W17(W17TO59), .W18(W18TO59), .W19(W19TO59), .W20(W20TO59), .W21(W21TO59), .W22(W22TO59), .W23(W23TO59), .W24(W24TO59), .W25(W25TO59), .W26(W26TO59), .W27(W27TO59), .W28(W28TO59), .W29(W29TO59), .W30(W30TO59), .W31(W31TO59), .W32(W32TO59), .W33(W33TO59), .W34(W34TO59), .W35(W35TO59), .W36(W36TO59), .W37(W37TO59), .W38(W38TO59), .W39(W39TO59), .W40(W40TO59), .W41(W41TO59), .W42(W42TO59), .W43(W43TO59), .W44(W44TO59), .W45(W45TO59), .W46(W46TO59), .W47(W47TO59), .W48(W48TO59), .W49(W49TO59), .W50(W50TO59), .W51(W51TO59), .W52(W52TO59), .W53(W53TO59), .W54(W54TO59), .W55(W55TO59), .W56(W56TO59), .W57(W57TO59), .W58(W58TO59), .W59(W59TO59), .W60(W60TO59), .W61(W61TO59), .W62(W62TO59), .W63(W63TO59)) neuron59(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out59));
neuron64in #(.W0(W0TO60), .W1(W1TO60), .W2(W2TO60), .W3(W3TO60), .W4(W4TO60), .W5(W5TO60), .W6(W6TO60), .W7(W7TO60), .W8(W8TO60), .W9(W9TO60), .W10(W10TO60), .W11(W11TO60), .W12(W12TO60), .W13(W13TO60), .W14(W14TO60), .W15(W15TO60), .W16(W16TO60), .W17(W17TO60), .W18(W18TO60), .W19(W19TO60), .W20(W20TO60), .W21(W21TO60), .W22(W22TO60), .W23(W23TO60), .W24(W24TO60), .W25(W25TO60), .W26(W26TO60), .W27(W27TO60), .W28(W28TO60), .W29(W29TO60), .W30(W30TO60), .W31(W31TO60), .W32(W32TO60), .W33(W33TO60), .W34(W34TO60), .W35(W35TO60), .W36(W36TO60), .W37(W37TO60), .W38(W38TO60), .W39(W39TO60), .W40(W40TO60), .W41(W41TO60), .W42(W42TO60), .W43(W43TO60), .W44(W44TO60), .W45(W45TO60), .W46(W46TO60), .W47(W47TO60), .W48(W48TO60), .W49(W49TO60), .W50(W50TO60), .W51(W51TO60), .W52(W52TO60), .W53(W53TO60), .W54(W54TO60), .W55(W55TO60), .W56(W56TO60), .W57(W57TO60), .W58(W58TO60), .W59(W59TO60), .W60(W60TO60), .W61(W61TO60), .W62(W62TO60), .W63(W63TO60)) neuron60(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out60));
neuron64in #(.W0(W0TO61), .W1(W1TO61), .W2(W2TO61), .W3(W3TO61), .W4(W4TO61), .W5(W5TO61), .W6(W6TO61), .W7(W7TO61), .W8(W8TO61), .W9(W9TO61), .W10(W10TO61), .W11(W11TO61), .W12(W12TO61), .W13(W13TO61), .W14(W14TO61), .W15(W15TO61), .W16(W16TO61), .W17(W17TO61), .W18(W18TO61), .W19(W19TO61), .W20(W20TO61), .W21(W21TO61), .W22(W22TO61), .W23(W23TO61), .W24(W24TO61), .W25(W25TO61), .W26(W26TO61), .W27(W27TO61), .W28(W28TO61), .W29(W29TO61), .W30(W30TO61), .W31(W31TO61), .W32(W32TO61), .W33(W33TO61), .W34(W34TO61), .W35(W35TO61), .W36(W36TO61), .W37(W37TO61), .W38(W38TO61), .W39(W39TO61), .W40(W40TO61), .W41(W41TO61), .W42(W42TO61), .W43(W43TO61), .W44(W44TO61), .W45(W45TO61), .W46(W46TO61), .W47(W47TO61), .W48(W48TO61), .W49(W49TO61), .W50(W50TO61), .W51(W51TO61), .W52(W52TO61), .W53(W53TO61), .W54(W54TO61), .W55(W55TO61), .W56(W56TO61), .W57(W57TO61), .W58(W58TO61), .W59(W59TO61), .W60(W60TO61), .W61(W61TO61), .W62(W62TO61), .W63(W63TO61)) neuron61(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out61));
neuron64in #(.W0(W0TO62), .W1(W1TO62), .W2(W2TO62), .W3(W3TO62), .W4(W4TO62), .W5(W5TO62), .W6(W6TO62), .W7(W7TO62), .W8(W8TO62), .W9(W9TO62), .W10(W10TO62), .W11(W11TO62), .W12(W12TO62), .W13(W13TO62), .W14(W14TO62), .W15(W15TO62), .W16(W16TO62), .W17(W17TO62), .W18(W18TO62), .W19(W19TO62), .W20(W20TO62), .W21(W21TO62), .W22(W22TO62), .W23(W23TO62), .W24(W24TO62), .W25(W25TO62), .W26(W26TO62), .W27(W27TO62), .W28(W28TO62), .W29(W29TO62), .W30(W30TO62), .W31(W31TO62), .W32(W32TO62), .W33(W33TO62), .W34(W34TO62), .W35(W35TO62), .W36(W36TO62), .W37(W37TO62), .W38(W38TO62), .W39(W39TO62), .W40(W40TO62), .W41(W41TO62), .W42(W42TO62), .W43(W43TO62), .W44(W44TO62), .W45(W45TO62), .W46(W46TO62), .W47(W47TO62), .W48(W48TO62), .W49(W49TO62), .W50(W50TO62), .W51(W51TO62), .W52(W52TO62), .W53(W53TO62), .W54(W54TO62), .W55(W55TO62), .W56(W56TO62), .W57(W57TO62), .W58(W58TO62), .W59(W59TO62), .W60(W60TO62), .W61(W61TO62), .W62(W62TO62), .W63(W63TO62)) neuron62(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out62));
neuron64in #(.W0(W0TO63), .W1(W1TO63), .W2(W2TO63), .W3(W3TO63), .W4(W4TO63), .W5(W5TO63), .W6(W6TO63), .W7(W7TO63), .W8(W8TO63), .W9(W9TO63), .W10(W10TO63), .W11(W11TO63), .W12(W12TO63), .W13(W13TO63), .W14(W14TO63), .W15(W15TO63), .W16(W16TO63), .W17(W17TO63), .W18(W18TO63), .W19(W19TO63), .W20(W20TO63), .W21(W21TO63), .W22(W22TO63), .W23(W23TO63), .W24(W24TO63), .W25(W25TO63), .W26(W26TO63), .W27(W27TO63), .W28(W28TO63), .W29(W29TO63), .W30(W30TO63), .W31(W31TO63), .W32(W32TO63), .W33(W33TO63), .W34(W34TO63), .W35(W35TO63), .W36(W36TO63), .W37(W37TO63), .W38(W38TO63), .W39(W39TO63), .W40(W40TO63), .W41(W41TO63), .W42(W42TO63), .W43(W43TO63), .W44(W44TO63), .W45(W45TO63), .W46(W46TO63), .W47(W47TO63), .W48(W48TO63), .W49(W49TO63), .W50(W50TO63), .W51(W51TO63), .W52(W52TO63), .W53(W53TO63), .W54(W54TO63), .W55(W55TO63), .W56(W56TO63), .W57(W57TO63), .W58(W58TO63), .W59(W59TO63), .W60(W60TO63), .W61(W61TO63), .W62(W62TO63), .W63(W63TO63)) neuron63(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out63));
neuron64in #(.W0(W0TO64), .W1(W1TO64), .W2(W2TO64), .W3(W3TO64), .W4(W4TO64), .W5(W5TO64), .W6(W6TO64), .W7(W7TO64), .W8(W8TO64), .W9(W9TO64), .W10(W10TO64), .W11(W11TO64), .W12(W12TO64), .W13(W13TO64), .W14(W14TO64), .W15(W15TO64), .W16(W16TO64), .W17(W17TO64), .W18(W18TO64), .W19(W19TO64), .W20(W20TO64), .W21(W21TO64), .W22(W22TO64), .W23(W23TO64), .W24(W24TO64), .W25(W25TO64), .W26(W26TO64), .W27(W27TO64), .W28(W28TO64), .W29(W29TO64), .W30(W30TO64), .W31(W31TO64), .W32(W32TO64), .W33(W33TO64), .W34(W34TO64), .W35(W35TO64), .W36(W36TO64), .W37(W37TO64), .W38(W38TO64), .W39(W39TO64), .W40(W40TO64), .W41(W41TO64), .W42(W42TO64), .W43(W43TO64), .W44(W44TO64), .W45(W45TO64), .W46(W46TO64), .W47(W47TO64), .W48(W48TO64), .W49(W49TO64), .W50(W50TO64), .W51(W51TO64), .W52(W52TO64), .W53(W53TO64), .W54(W54TO64), .W55(W55TO64), .W56(W56TO64), .W57(W57TO64), .W58(W58TO64), .W59(W59TO64), .W60(W60TO64), .W61(W61TO64), .W62(W62TO64), .W63(W63TO64)) neuron64(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out64));
neuron64in #(.W0(W0TO65), .W1(W1TO65), .W2(W2TO65), .W3(W3TO65), .W4(W4TO65), .W5(W5TO65), .W6(W6TO65), .W7(W7TO65), .W8(W8TO65), .W9(W9TO65), .W10(W10TO65), .W11(W11TO65), .W12(W12TO65), .W13(W13TO65), .W14(W14TO65), .W15(W15TO65), .W16(W16TO65), .W17(W17TO65), .W18(W18TO65), .W19(W19TO65), .W20(W20TO65), .W21(W21TO65), .W22(W22TO65), .W23(W23TO65), .W24(W24TO65), .W25(W25TO65), .W26(W26TO65), .W27(W27TO65), .W28(W28TO65), .W29(W29TO65), .W30(W30TO65), .W31(W31TO65), .W32(W32TO65), .W33(W33TO65), .W34(W34TO65), .W35(W35TO65), .W36(W36TO65), .W37(W37TO65), .W38(W38TO65), .W39(W39TO65), .W40(W40TO65), .W41(W41TO65), .W42(W42TO65), .W43(W43TO65), .W44(W44TO65), .W45(W45TO65), .W46(W46TO65), .W47(W47TO65), .W48(W48TO65), .W49(W49TO65), .W50(W50TO65), .W51(W51TO65), .W52(W52TO65), .W53(W53TO65), .W54(W54TO65), .W55(W55TO65), .W56(W56TO65), .W57(W57TO65), .W58(W58TO65), .W59(W59TO65), .W60(W60TO65), .W61(W61TO65), .W62(W62TO65), .W63(W63TO65)) neuron65(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out65));
neuron64in #(.W0(W0TO66), .W1(W1TO66), .W2(W2TO66), .W3(W3TO66), .W4(W4TO66), .W5(W5TO66), .W6(W6TO66), .W7(W7TO66), .W8(W8TO66), .W9(W9TO66), .W10(W10TO66), .W11(W11TO66), .W12(W12TO66), .W13(W13TO66), .W14(W14TO66), .W15(W15TO66), .W16(W16TO66), .W17(W17TO66), .W18(W18TO66), .W19(W19TO66), .W20(W20TO66), .W21(W21TO66), .W22(W22TO66), .W23(W23TO66), .W24(W24TO66), .W25(W25TO66), .W26(W26TO66), .W27(W27TO66), .W28(W28TO66), .W29(W29TO66), .W30(W30TO66), .W31(W31TO66), .W32(W32TO66), .W33(W33TO66), .W34(W34TO66), .W35(W35TO66), .W36(W36TO66), .W37(W37TO66), .W38(W38TO66), .W39(W39TO66), .W40(W40TO66), .W41(W41TO66), .W42(W42TO66), .W43(W43TO66), .W44(W44TO66), .W45(W45TO66), .W46(W46TO66), .W47(W47TO66), .W48(W48TO66), .W49(W49TO66), .W50(W50TO66), .W51(W51TO66), .W52(W52TO66), .W53(W53TO66), .W54(W54TO66), .W55(W55TO66), .W56(W56TO66), .W57(W57TO66), .W58(W58TO66), .W59(W59TO66), .W60(W60TO66), .W61(W61TO66), .W62(W62TO66), .W63(W63TO66)) neuron66(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out66));
neuron64in #(.W0(W0TO67), .W1(W1TO67), .W2(W2TO67), .W3(W3TO67), .W4(W4TO67), .W5(W5TO67), .W6(W6TO67), .W7(W7TO67), .W8(W8TO67), .W9(W9TO67), .W10(W10TO67), .W11(W11TO67), .W12(W12TO67), .W13(W13TO67), .W14(W14TO67), .W15(W15TO67), .W16(W16TO67), .W17(W17TO67), .W18(W18TO67), .W19(W19TO67), .W20(W20TO67), .W21(W21TO67), .W22(W22TO67), .W23(W23TO67), .W24(W24TO67), .W25(W25TO67), .W26(W26TO67), .W27(W27TO67), .W28(W28TO67), .W29(W29TO67), .W30(W30TO67), .W31(W31TO67), .W32(W32TO67), .W33(W33TO67), .W34(W34TO67), .W35(W35TO67), .W36(W36TO67), .W37(W37TO67), .W38(W38TO67), .W39(W39TO67), .W40(W40TO67), .W41(W41TO67), .W42(W42TO67), .W43(W43TO67), .W44(W44TO67), .W45(W45TO67), .W46(W46TO67), .W47(W47TO67), .W48(W48TO67), .W49(W49TO67), .W50(W50TO67), .W51(W51TO67), .W52(W52TO67), .W53(W53TO67), .W54(W54TO67), .W55(W55TO67), .W56(W56TO67), .W57(W57TO67), .W58(W58TO67), .W59(W59TO67), .W60(W60TO67), .W61(W61TO67), .W62(W62TO67), .W63(W63TO67)) neuron67(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out67));
neuron64in #(.W0(W0TO68), .W1(W1TO68), .W2(W2TO68), .W3(W3TO68), .W4(W4TO68), .W5(W5TO68), .W6(W6TO68), .W7(W7TO68), .W8(W8TO68), .W9(W9TO68), .W10(W10TO68), .W11(W11TO68), .W12(W12TO68), .W13(W13TO68), .W14(W14TO68), .W15(W15TO68), .W16(W16TO68), .W17(W17TO68), .W18(W18TO68), .W19(W19TO68), .W20(W20TO68), .W21(W21TO68), .W22(W22TO68), .W23(W23TO68), .W24(W24TO68), .W25(W25TO68), .W26(W26TO68), .W27(W27TO68), .W28(W28TO68), .W29(W29TO68), .W30(W30TO68), .W31(W31TO68), .W32(W32TO68), .W33(W33TO68), .W34(W34TO68), .W35(W35TO68), .W36(W36TO68), .W37(W37TO68), .W38(W38TO68), .W39(W39TO68), .W40(W40TO68), .W41(W41TO68), .W42(W42TO68), .W43(W43TO68), .W44(W44TO68), .W45(W45TO68), .W46(W46TO68), .W47(W47TO68), .W48(W48TO68), .W49(W49TO68), .W50(W50TO68), .W51(W51TO68), .W52(W52TO68), .W53(W53TO68), .W54(W54TO68), .W55(W55TO68), .W56(W56TO68), .W57(W57TO68), .W58(W58TO68), .W59(W59TO68), .W60(W60TO68), .W61(W61TO68), .W62(W62TO68), .W63(W63TO68)) neuron68(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out68));
neuron64in #(.W0(W0TO69), .W1(W1TO69), .W2(W2TO69), .W3(W3TO69), .W4(W4TO69), .W5(W5TO69), .W6(W6TO69), .W7(W7TO69), .W8(W8TO69), .W9(W9TO69), .W10(W10TO69), .W11(W11TO69), .W12(W12TO69), .W13(W13TO69), .W14(W14TO69), .W15(W15TO69), .W16(W16TO69), .W17(W17TO69), .W18(W18TO69), .W19(W19TO69), .W20(W20TO69), .W21(W21TO69), .W22(W22TO69), .W23(W23TO69), .W24(W24TO69), .W25(W25TO69), .W26(W26TO69), .W27(W27TO69), .W28(W28TO69), .W29(W29TO69), .W30(W30TO69), .W31(W31TO69), .W32(W32TO69), .W33(W33TO69), .W34(W34TO69), .W35(W35TO69), .W36(W36TO69), .W37(W37TO69), .W38(W38TO69), .W39(W39TO69), .W40(W40TO69), .W41(W41TO69), .W42(W42TO69), .W43(W43TO69), .W44(W44TO69), .W45(W45TO69), .W46(W46TO69), .W47(W47TO69), .W48(W48TO69), .W49(W49TO69), .W50(W50TO69), .W51(W51TO69), .W52(W52TO69), .W53(W53TO69), .W54(W54TO69), .W55(W55TO69), .W56(W56TO69), .W57(W57TO69), .W58(W58TO69), .W59(W59TO69), .W60(W60TO69), .W61(W61TO69), .W62(W62TO69), .W63(W63TO69)) neuron69(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out69));
neuron64in #(.W0(W0TO70), .W1(W1TO70), .W2(W2TO70), .W3(W3TO70), .W4(W4TO70), .W5(W5TO70), .W6(W6TO70), .W7(W7TO70), .W8(W8TO70), .W9(W9TO70), .W10(W10TO70), .W11(W11TO70), .W12(W12TO70), .W13(W13TO70), .W14(W14TO70), .W15(W15TO70), .W16(W16TO70), .W17(W17TO70), .W18(W18TO70), .W19(W19TO70), .W20(W20TO70), .W21(W21TO70), .W22(W22TO70), .W23(W23TO70), .W24(W24TO70), .W25(W25TO70), .W26(W26TO70), .W27(W27TO70), .W28(W28TO70), .W29(W29TO70), .W30(W30TO70), .W31(W31TO70), .W32(W32TO70), .W33(W33TO70), .W34(W34TO70), .W35(W35TO70), .W36(W36TO70), .W37(W37TO70), .W38(W38TO70), .W39(W39TO70), .W40(W40TO70), .W41(W41TO70), .W42(W42TO70), .W43(W43TO70), .W44(W44TO70), .W45(W45TO70), .W46(W46TO70), .W47(W47TO70), .W48(W48TO70), .W49(W49TO70), .W50(W50TO70), .W51(W51TO70), .W52(W52TO70), .W53(W53TO70), .W54(W54TO70), .W55(W55TO70), .W56(W56TO70), .W57(W57TO70), .W58(W58TO70), .W59(W59TO70), .W60(W60TO70), .W61(W61TO70), .W62(W62TO70), .W63(W63TO70)) neuron70(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out70));
neuron64in #(.W0(W0TO71), .W1(W1TO71), .W2(W2TO71), .W3(W3TO71), .W4(W4TO71), .W5(W5TO71), .W6(W6TO71), .W7(W7TO71), .W8(W8TO71), .W9(W9TO71), .W10(W10TO71), .W11(W11TO71), .W12(W12TO71), .W13(W13TO71), .W14(W14TO71), .W15(W15TO71), .W16(W16TO71), .W17(W17TO71), .W18(W18TO71), .W19(W19TO71), .W20(W20TO71), .W21(W21TO71), .W22(W22TO71), .W23(W23TO71), .W24(W24TO71), .W25(W25TO71), .W26(W26TO71), .W27(W27TO71), .W28(W28TO71), .W29(W29TO71), .W30(W30TO71), .W31(W31TO71), .W32(W32TO71), .W33(W33TO71), .W34(W34TO71), .W35(W35TO71), .W36(W36TO71), .W37(W37TO71), .W38(W38TO71), .W39(W39TO71), .W40(W40TO71), .W41(W41TO71), .W42(W42TO71), .W43(W43TO71), .W44(W44TO71), .W45(W45TO71), .W46(W46TO71), .W47(W47TO71), .W48(W48TO71), .W49(W49TO71), .W50(W50TO71), .W51(W51TO71), .W52(W52TO71), .W53(W53TO71), .W54(W54TO71), .W55(W55TO71), .W56(W56TO71), .W57(W57TO71), .W58(W58TO71), .W59(W59TO71), .W60(W60TO71), .W61(W61TO71), .W62(W62TO71), .W63(W63TO71)) neuron71(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out71));
neuron64in #(.W0(W0TO72), .W1(W1TO72), .W2(W2TO72), .W3(W3TO72), .W4(W4TO72), .W5(W5TO72), .W6(W6TO72), .W7(W7TO72), .W8(W8TO72), .W9(W9TO72), .W10(W10TO72), .W11(W11TO72), .W12(W12TO72), .W13(W13TO72), .W14(W14TO72), .W15(W15TO72), .W16(W16TO72), .W17(W17TO72), .W18(W18TO72), .W19(W19TO72), .W20(W20TO72), .W21(W21TO72), .W22(W22TO72), .W23(W23TO72), .W24(W24TO72), .W25(W25TO72), .W26(W26TO72), .W27(W27TO72), .W28(W28TO72), .W29(W29TO72), .W30(W30TO72), .W31(W31TO72), .W32(W32TO72), .W33(W33TO72), .W34(W34TO72), .W35(W35TO72), .W36(W36TO72), .W37(W37TO72), .W38(W38TO72), .W39(W39TO72), .W40(W40TO72), .W41(W41TO72), .W42(W42TO72), .W43(W43TO72), .W44(W44TO72), .W45(W45TO72), .W46(W46TO72), .W47(W47TO72), .W48(W48TO72), .W49(W49TO72), .W50(W50TO72), .W51(W51TO72), .W52(W52TO72), .W53(W53TO72), .W54(W54TO72), .W55(W55TO72), .W56(W56TO72), .W57(W57TO72), .W58(W58TO72), .W59(W59TO72), .W60(W60TO72), .W61(W61TO72), .W62(W62TO72), .W63(W63TO72)) neuron72(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out72));
neuron64in #(.W0(W0TO73), .W1(W1TO73), .W2(W2TO73), .W3(W3TO73), .W4(W4TO73), .W5(W5TO73), .W6(W6TO73), .W7(W7TO73), .W8(W8TO73), .W9(W9TO73), .W10(W10TO73), .W11(W11TO73), .W12(W12TO73), .W13(W13TO73), .W14(W14TO73), .W15(W15TO73), .W16(W16TO73), .W17(W17TO73), .W18(W18TO73), .W19(W19TO73), .W20(W20TO73), .W21(W21TO73), .W22(W22TO73), .W23(W23TO73), .W24(W24TO73), .W25(W25TO73), .W26(W26TO73), .W27(W27TO73), .W28(W28TO73), .W29(W29TO73), .W30(W30TO73), .W31(W31TO73), .W32(W32TO73), .W33(W33TO73), .W34(W34TO73), .W35(W35TO73), .W36(W36TO73), .W37(W37TO73), .W38(W38TO73), .W39(W39TO73), .W40(W40TO73), .W41(W41TO73), .W42(W42TO73), .W43(W43TO73), .W44(W44TO73), .W45(W45TO73), .W46(W46TO73), .W47(W47TO73), .W48(W48TO73), .W49(W49TO73), .W50(W50TO73), .W51(W51TO73), .W52(W52TO73), .W53(W53TO73), .W54(W54TO73), .W55(W55TO73), .W56(W56TO73), .W57(W57TO73), .W58(W58TO73), .W59(W59TO73), .W60(W60TO73), .W61(W61TO73), .W62(W62TO73), .W63(W63TO73)) neuron73(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out73));
neuron64in #(.W0(W0TO74), .W1(W1TO74), .W2(W2TO74), .W3(W3TO74), .W4(W4TO74), .W5(W5TO74), .W6(W6TO74), .W7(W7TO74), .W8(W8TO74), .W9(W9TO74), .W10(W10TO74), .W11(W11TO74), .W12(W12TO74), .W13(W13TO74), .W14(W14TO74), .W15(W15TO74), .W16(W16TO74), .W17(W17TO74), .W18(W18TO74), .W19(W19TO74), .W20(W20TO74), .W21(W21TO74), .W22(W22TO74), .W23(W23TO74), .W24(W24TO74), .W25(W25TO74), .W26(W26TO74), .W27(W27TO74), .W28(W28TO74), .W29(W29TO74), .W30(W30TO74), .W31(W31TO74), .W32(W32TO74), .W33(W33TO74), .W34(W34TO74), .W35(W35TO74), .W36(W36TO74), .W37(W37TO74), .W38(W38TO74), .W39(W39TO74), .W40(W40TO74), .W41(W41TO74), .W42(W42TO74), .W43(W43TO74), .W44(W44TO74), .W45(W45TO74), .W46(W46TO74), .W47(W47TO74), .W48(W48TO74), .W49(W49TO74), .W50(W50TO74), .W51(W51TO74), .W52(W52TO74), .W53(W53TO74), .W54(W54TO74), .W55(W55TO74), .W56(W56TO74), .W57(W57TO74), .W58(W58TO74), .W59(W59TO74), .W60(W60TO74), .W61(W61TO74), .W62(W62TO74), .W63(W63TO74)) neuron74(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out74));
neuron64in #(.W0(W0TO75), .W1(W1TO75), .W2(W2TO75), .W3(W3TO75), .W4(W4TO75), .W5(W5TO75), .W6(W6TO75), .W7(W7TO75), .W8(W8TO75), .W9(W9TO75), .W10(W10TO75), .W11(W11TO75), .W12(W12TO75), .W13(W13TO75), .W14(W14TO75), .W15(W15TO75), .W16(W16TO75), .W17(W17TO75), .W18(W18TO75), .W19(W19TO75), .W20(W20TO75), .W21(W21TO75), .W22(W22TO75), .W23(W23TO75), .W24(W24TO75), .W25(W25TO75), .W26(W26TO75), .W27(W27TO75), .W28(W28TO75), .W29(W29TO75), .W30(W30TO75), .W31(W31TO75), .W32(W32TO75), .W33(W33TO75), .W34(W34TO75), .W35(W35TO75), .W36(W36TO75), .W37(W37TO75), .W38(W38TO75), .W39(W39TO75), .W40(W40TO75), .W41(W41TO75), .W42(W42TO75), .W43(W43TO75), .W44(W44TO75), .W45(W45TO75), .W46(W46TO75), .W47(W47TO75), .W48(W48TO75), .W49(W49TO75), .W50(W50TO75), .W51(W51TO75), .W52(W52TO75), .W53(W53TO75), .W54(W54TO75), .W55(W55TO75), .W56(W56TO75), .W57(W57TO75), .W58(W58TO75), .W59(W59TO75), .W60(W60TO75), .W61(W61TO75), .W62(W62TO75), .W63(W63TO75)) neuron75(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out75));
neuron64in #(.W0(W0TO76), .W1(W1TO76), .W2(W2TO76), .W3(W3TO76), .W4(W4TO76), .W5(W5TO76), .W6(W6TO76), .W7(W7TO76), .W8(W8TO76), .W9(W9TO76), .W10(W10TO76), .W11(W11TO76), .W12(W12TO76), .W13(W13TO76), .W14(W14TO76), .W15(W15TO76), .W16(W16TO76), .W17(W17TO76), .W18(W18TO76), .W19(W19TO76), .W20(W20TO76), .W21(W21TO76), .W22(W22TO76), .W23(W23TO76), .W24(W24TO76), .W25(W25TO76), .W26(W26TO76), .W27(W27TO76), .W28(W28TO76), .W29(W29TO76), .W30(W30TO76), .W31(W31TO76), .W32(W32TO76), .W33(W33TO76), .W34(W34TO76), .W35(W35TO76), .W36(W36TO76), .W37(W37TO76), .W38(W38TO76), .W39(W39TO76), .W40(W40TO76), .W41(W41TO76), .W42(W42TO76), .W43(W43TO76), .W44(W44TO76), .W45(W45TO76), .W46(W46TO76), .W47(W47TO76), .W48(W48TO76), .W49(W49TO76), .W50(W50TO76), .W51(W51TO76), .W52(W52TO76), .W53(W53TO76), .W54(W54TO76), .W55(W55TO76), .W56(W56TO76), .W57(W57TO76), .W58(W58TO76), .W59(W59TO76), .W60(W60TO76), .W61(W61TO76), .W62(W62TO76), .W63(W63TO76)) neuron76(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out76));
neuron64in #(.W0(W0TO77), .W1(W1TO77), .W2(W2TO77), .W3(W3TO77), .W4(W4TO77), .W5(W5TO77), .W6(W6TO77), .W7(W7TO77), .W8(W8TO77), .W9(W9TO77), .W10(W10TO77), .W11(W11TO77), .W12(W12TO77), .W13(W13TO77), .W14(W14TO77), .W15(W15TO77), .W16(W16TO77), .W17(W17TO77), .W18(W18TO77), .W19(W19TO77), .W20(W20TO77), .W21(W21TO77), .W22(W22TO77), .W23(W23TO77), .W24(W24TO77), .W25(W25TO77), .W26(W26TO77), .W27(W27TO77), .W28(W28TO77), .W29(W29TO77), .W30(W30TO77), .W31(W31TO77), .W32(W32TO77), .W33(W33TO77), .W34(W34TO77), .W35(W35TO77), .W36(W36TO77), .W37(W37TO77), .W38(W38TO77), .W39(W39TO77), .W40(W40TO77), .W41(W41TO77), .W42(W42TO77), .W43(W43TO77), .W44(W44TO77), .W45(W45TO77), .W46(W46TO77), .W47(W47TO77), .W48(W48TO77), .W49(W49TO77), .W50(W50TO77), .W51(W51TO77), .W52(W52TO77), .W53(W53TO77), .W54(W54TO77), .W55(W55TO77), .W56(W56TO77), .W57(W57TO77), .W58(W58TO77), .W59(W59TO77), .W60(W60TO77), .W61(W61TO77), .W62(W62TO77), .W63(W63TO77)) neuron77(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out77));
neuron64in #(.W0(W0TO78), .W1(W1TO78), .W2(W2TO78), .W3(W3TO78), .W4(W4TO78), .W5(W5TO78), .W6(W6TO78), .W7(W7TO78), .W8(W8TO78), .W9(W9TO78), .W10(W10TO78), .W11(W11TO78), .W12(W12TO78), .W13(W13TO78), .W14(W14TO78), .W15(W15TO78), .W16(W16TO78), .W17(W17TO78), .W18(W18TO78), .W19(W19TO78), .W20(W20TO78), .W21(W21TO78), .W22(W22TO78), .W23(W23TO78), .W24(W24TO78), .W25(W25TO78), .W26(W26TO78), .W27(W27TO78), .W28(W28TO78), .W29(W29TO78), .W30(W30TO78), .W31(W31TO78), .W32(W32TO78), .W33(W33TO78), .W34(W34TO78), .W35(W35TO78), .W36(W36TO78), .W37(W37TO78), .W38(W38TO78), .W39(W39TO78), .W40(W40TO78), .W41(W41TO78), .W42(W42TO78), .W43(W43TO78), .W44(W44TO78), .W45(W45TO78), .W46(W46TO78), .W47(W47TO78), .W48(W48TO78), .W49(W49TO78), .W50(W50TO78), .W51(W51TO78), .W52(W52TO78), .W53(W53TO78), .W54(W54TO78), .W55(W55TO78), .W56(W56TO78), .W57(W57TO78), .W58(W58TO78), .W59(W59TO78), .W60(W60TO78), .W61(W61TO78), .W62(W62TO78), .W63(W63TO78)) neuron78(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out78));
neuron64in #(.W0(W0TO79), .W1(W1TO79), .W2(W2TO79), .W3(W3TO79), .W4(W4TO79), .W5(W5TO79), .W6(W6TO79), .W7(W7TO79), .W8(W8TO79), .W9(W9TO79), .W10(W10TO79), .W11(W11TO79), .W12(W12TO79), .W13(W13TO79), .W14(W14TO79), .W15(W15TO79), .W16(W16TO79), .W17(W17TO79), .W18(W18TO79), .W19(W19TO79), .W20(W20TO79), .W21(W21TO79), .W22(W22TO79), .W23(W23TO79), .W24(W24TO79), .W25(W25TO79), .W26(W26TO79), .W27(W27TO79), .W28(W28TO79), .W29(W29TO79), .W30(W30TO79), .W31(W31TO79), .W32(W32TO79), .W33(W33TO79), .W34(W34TO79), .W35(W35TO79), .W36(W36TO79), .W37(W37TO79), .W38(W38TO79), .W39(W39TO79), .W40(W40TO79), .W41(W41TO79), .W42(W42TO79), .W43(W43TO79), .W44(W44TO79), .W45(W45TO79), .W46(W46TO79), .W47(W47TO79), .W48(W48TO79), .W49(W49TO79), .W50(W50TO79), .W51(W51TO79), .W52(W52TO79), .W53(W53TO79), .W54(W54TO79), .W55(W55TO79), .W56(W56TO79), .W57(W57TO79), .W58(W58TO79), .W59(W59TO79), .W60(W60TO79), .W61(W61TO79), .W62(W62TO79), .W63(W63TO79)) neuron79(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out79));
neuron64in #(.W0(W0TO80), .W1(W1TO80), .W2(W2TO80), .W3(W3TO80), .W4(W4TO80), .W5(W5TO80), .W6(W6TO80), .W7(W7TO80), .W8(W8TO80), .W9(W9TO80), .W10(W10TO80), .W11(W11TO80), .W12(W12TO80), .W13(W13TO80), .W14(W14TO80), .W15(W15TO80), .W16(W16TO80), .W17(W17TO80), .W18(W18TO80), .W19(W19TO80), .W20(W20TO80), .W21(W21TO80), .W22(W22TO80), .W23(W23TO80), .W24(W24TO80), .W25(W25TO80), .W26(W26TO80), .W27(W27TO80), .W28(W28TO80), .W29(W29TO80), .W30(W30TO80), .W31(W31TO80), .W32(W32TO80), .W33(W33TO80), .W34(W34TO80), .W35(W35TO80), .W36(W36TO80), .W37(W37TO80), .W38(W38TO80), .W39(W39TO80), .W40(W40TO80), .W41(W41TO80), .W42(W42TO80), .W43(W43TO80), .W44(W44TO80), .W45(W45TO80), .W46(W46TO80), .W47(W47TO80), .W48(W48TO80), .W49(W49TO80), .W50(W50TO80), .W51(W51TO80), .W52(W52TO80), .W53(W53TO80), .W54(W54TO80), .W55(W55TO80), .W56(W56TO80), .W57(W57TO80), .W58(W58TO80), .W59(W59TO80), .W60(W60TO80), .W61(W61TO80), .W62(W62TO80), .W63(W63TO80)) neuron80(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out80));
neuron64in #(.W0(W0TO81), .W1(W1TO81), .W2(W2TO81), .W3(W3TO81), .W4(W4TO81), .W5(W5TO81), .W6(W6TO81), .W7(W7TO81), .W8(W8TO81), .W9(W9TO81), .W10(W10TO81), .W11(W11TO81), .W12(W12TO81), .W13(W13TO81), .W14(W14TO81), .W15(W15TO81), .W16(W16TO81), .W17(W17TO81), .W18(W18TO81), .W19(W19TO81), .W20(W20TO81), .W21(W21TO81), .W22(W22TO81), .W23(W23TO81), .W24(W24TO81), .W25(W25TO81), .W26(W26TO81), .W27(W27TO81), .W28(W28TO81), .W29(W29TO81), .W30(W30TO81), .W31(W31TO81), .W32(W32TO81), .W33(W33TO81), .W34(W34TO81), .W35(W35TO81), .W36(W36TO81), .W37(W37TO81), .W38(W38TO81), .W39(W39TO81), .W40(W40TO81), .W41(W41TO81), .W42(W42TO81), .W43(W43TO81), .W44(W44TO81), .W45(W45TO81), .W46(W46TO81), .W47(W47TO81), .W48(W48TO81), .W49(W49TO81), .W50(W50TO81), .W51(W51TO81), .W52(W52TO81), .W53(W53TO81), .W54(W54TO81), .W55(W55TO81), .W56(W56TO81), .W57(W57TO81), .W58(W58TO81), .W59(W59TO81), .W60(W60TO81), .W61(W61TO81), .W62(W62TO81), .W63(W63TO81)) neuron81(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out81));
neuron64in #(.W0(W0TO82), .W1(W1TO82), .W2(W2TO82), .W3(W3TO82), .W4(W4TO82), .W5(W5TO82), .W6(W6TO82), .W7(W7TO82), .W8(W8TO82), .W9(W9TO82), .W10(W10TO82), .W11(W11TO82), .W12(W12TO82), .W13(W13TO82), .W14(W14TO82), .W15(W15TO82), .W16(W16TO82), .W17(W17TO82), .W18(W18TO82), .W19(W19TO82), .W20(W20TO82), .W21(W21TO82), .W22(W22TO82), .W23(W23TO82), .W24(W24TO82), .W25(W25TO82), .W26(W26TO82), .W27(W27TO82), .W28(W28TO82), .W29(W29TO82), .W30(W30TO82), .W31(W31TO82), .W32(W32TO82), .W33(W33TO82), .W34(W34TO82), .W35(W35TO82), .W36(W36TO82), .W37(W37TO82), .W38(W38TO82), .W39(W39TO82), .W40(W40TO82), .W41(W41TO82), .W42(W42TO82), .W43(W43TO82), .W44(W44TO82), .W45(W45TO82), .W46(W46TO82), .W47(W47TO82), .W48(W48TO82), .W49(W49TO82), .W50(W50TO82), .W51(W51TO82), .W52(W52TO82), .W53(W53TO82), .W54(W54TO82), .W55(W55TO82), .W56(W56TO82), .W57(W57TO82), .W58(W58TO82), .W59(W59TO82), .W60(W60TO82), .W61(W61TO82), .W62(W62TO82), .W63(W63TO82)) neuron82(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out82));
neuron64in #(.W0(W0TO83), .W1(W1TO83), .W2(W2TO83), .W3(W3TO83), .W4(W4TO83), .W5(W5TO83), .W6(W6TO83), .W7(W7TO83), .W8(W8TO83), .W9(W9TO83), .W10(W10TO83), .W11(W11TO83), .W12(W12TO83), .W13(W13TO83), .W14(W14TO83), .W15(W15TO83), .W16(W16TO83), .W17(W17TO83), .W18(W18TO83), .W19(W19TO83), .W20(W20TO83), .W21(W21TO83), .W22(W22TO83), .W23(W23TO83), .W24(W24TO83), .W25(W25TO83), .W26(W26TO83), .W27(W27TO83), .W28(W28TO83), .W29(W29TO83), .W30(W30TO83), .W31(W31TO83), .W32(W32TO83), .W33(W33TO83), .W34(W34TO83), .W35(W35TO83), .W36(W36TO83), .W37(W37TO83), .W38(W38TO83), .W39(W39TO83), .W40(W40TO83), .W41(W41TO83), .W42(W42TO83), .W43(W43TO83), .W44(W44TO83), .W45(W45TO83), .W46(W46TO83), .W47(W47TO83), .W48(W48TO83), .W49(W49TO83), .W50(W50TO83), .W51(W51TO83), .W52(W52TO83), .W53(W53TO83), .W54(W54TO83), .W55(W55TO83), .W56(W56TO83), .W57(W57TO83), .W58(W58TO83), .W59(W59TO83), .W60(W60TO83), .W61(W61TO83), .W62(W62TO83), .W63(W63TO83)) neuron83(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out83));
neuron64in #(.W0(W0TO84), .W1(W1TO84), .W2(W2TO84), .W3(W3TO84), .W4(W4TO84), .W5(W5TO84), .W6(W6TO84), .W7(W7TO84), .W8(W8TO84), .W9(W9TO84), .W10(W10TO84), .W11(W11TO84), .W12(W12TO84), .W13(W13TO84), .W14(W14TO84), .W15(W15TO84), .W16(W16TO84), .W17(W17TO84), .W18(W18TO84), .W19(W19TO84), .W20(W20TO84), .W21(W21TO84), .W22(W22TO84), .W23(W23TO84), .W24(W24TO84), .W25(W25TO84), .W26(W26TO84), .W27(W27TO84), .W28(W28TO84), .W29(W29TO84), .W30(W30TO84), .W31(W31TO84), .W32(W32TO84), .W33(W33TO84), .W34(W34TO84), .W35(W35TO84), .W36(W36TO84), .W37(W37TO84), .W38(W38TO84), .W39(W39TO84), .W40(W40TO84), .W41(W41TO84), .W42(W42TO84), .W43(W43TO84), .W44(W44TO84), .W45(W45TO84), .W46(W46TO84), .W47(W47TO84), .W48(W48TO84), .W49(W49TO84), .W50(W50TO84), .W51(W51TO84), .W52(W52TO84), .W53(W53TO84), .W54(W54TO84), .W55(W55TO84), .W56(W56TO84), .W57(W57TO84), .W58(W58TO84), .W59(W59TO84), .W60(W60TO84), .W61(W61TO84), .W62(W62TO84), .W63(W63TO84)) neuron84(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out84));
neuron64in #(.W0(W0TO85), .W1(W1TO85), .W2(W2TO85), .W3(W3TO85), .W4(W4TO85), .W5(W5TO85), .W6(W6TO85), .W7(W7TO85), .W8(W8TO85), .W9(W9TO85), .W10(W10TO85), .W11(W11TO85), .W12(W12TO85), .W13(W13TO85), .W14(W14TO85), .W15(W15TO85), .W16(W16TO85), .W17(W17TO85), .W18(W18TO85), .W19(W19TO85), .W20(W20TO85), .W21(W21TO85), .W22(W22TO85), .W23(W23TO85), .W24(W24TO85), .W25(W25TO85), .W26(W26TO85), .W27(W27TO85), .W28(W28TO85), .W29(W29TO85), .W30(W30TO85), .W31(W31TO85), .W32(W32TO85), .W33(W33TO85), .W34(W34TO85), .W35(W35TO85), .W36(W36TO85), .W37(W37TO85), .W38(W38TO85), .W39(W39TO85), .W40(W40TO85), .W41(W41TO85), .W42(W42TO85), .W43(W43TO85), .W44(W44TO85), .W45(W45TO85), .W46(W46TO85), .W47(W47TO85), .W48(W48TO85), .W49(W49TO85), .W50(W50TO85), .W51(W51TO85), .W52(W52TO85), .W53(W53TO85), .W54(W54TO85), .W55(W55TO85), .W56(W56TO85), .W57(W57TO85), .W58(W58TO85), .W59(W59TO85), .W60(W60TO85), .W61(W61TO85), .W62(W62TO85), .W63(W63TO85)) neuron85(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out85));
neuron64in #(.W0(W0TO86), .W1(W1TO86), .W2(W2TO86), .W3(W3TO86), .W4(W4TO86), .W5(W5TO86), .W6(W6TO86), .W7(W7TO86), .W8(W8TO86), .W9(W9TO86), .W10(W10TO86), .W11(W11TO86), .W12(W12TO86), .W13(W13TO86), .W14(W14TO86), .W15(W15TO86), .W16(W16TO86), .W17(W17TO86), .W18(W18TO86), .W19(W19TO86), .W20(W20TO86), .W21(W21TO86), .W22(W22TO86), .W23(W23TO86), .W24(W24TO86), .W25(W25TO86), .W26(W26TO86), .W27(W27TO86), .W28(W28TO86), .W29(W29TO86), .W30(W30TO86), .W31(W31TO86), .W32(W32TO86), .W33(W33TO86), .W34(W34TO86), .W35(W35TO86), .W36(W36TO86), .W37(W37TO86), .W38(W38TO86), .W39(W39TO86), .W40(W40TO86), .W41(W41TO86), .W42(W42TO86), .W43(W43TO86), .W44(W44TO86), .W45(W45TO86), .W46(W46TO86), .W47(W47TO86), .W48(W48TO86), .W49(W49TO86), .W50(W50TO86), .W51(W51TO86), .W52(W52TO86), .W53(W53TO86), .W54(W54TO86), .W55(W55TO86), .W56(W56TO86), .W57(W57TO86), .W58(W58TO86), .W59(W59TO86), .W60(W60TO86), .W61(W61TO86), .W62(W62TO86), .W63(W63TO86)) neuron86(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out86));
neuron64in #(.W0(W0TO87), .W1(W1TO87), .W2(W2TO87), .W3(W3TO87), .W4(W4TO87), .W5(W5TO87), .W6(W6TO87), .W7(W7TO87), .W8(W8TO87), .W9(W9TO87), .W10(W10TO87), .W11(W11TO87), .W12(W12TO87), .W13(W13TO87), .W14(W14TO87), .W15(W15TO87), .W16(W16TO87), .W17(W17TO87), .W18(W18TO87), .W19(W19TO87), .W20(W20TO87), .W21(W21TO87), .W22(W22TO87), .W23(W23TO87), .W24(W24TO87), .W25(W25TO87), .W26(W26TO87), .W27(W27TO87), .W28(W28TO87), .W29(W29TO87), .W30(W30TO87), .W31(W31TO87), .W32(W32TO87), .W33(W33TO87), .W34(W34TO87), .W35(W35TO87), .W36(W36TO87), .W37(W37TO87), .W38(W38TO87), .W39(W39TO87), .W40(W40TO87), .W41(W41TO87), .W42(W42TO87), .W43(W43TO87), .W44(W44TO87), .W45(W45TO87), .W46(W46TO87), .W47(W47TO87), .W48(W48TO87), .W49(W49TO87), .W50(W50TO87), .W51(W51TO87), .W52(W52TO87), .W53(W53TO87), .W54(W54TO87), .W55(W55TO87), .W56(W56TO87), .W57(W57TO87), .W58(W58TO87), .W59(W59TO87), .W60(W60TO87), .W61(W61TO87), .W62(W62TO87), .W63(W63TO87)) neuron87(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out87));
neuron64in #(.W0(W0TO88), .W1(W1TO88), .W2(W2TO88), .W3(W3TO88), .W4(W4TO88), .W5(W5TO88), .W6(W6TO88), .W7(W7TO88), .W8(W8TO88), .W9(W9TO88), .W10(W10TO88), .W11(W11TO88), .W12(W12TO88), .W13(W13TO88), .W14(W14TO88), .W15(W15TO88), .W16(W16TO88), .W17(W17TO88), .W18(W18TO88), .W19(W19TO88), .W20(W20TO88), .W21(W21TO88), .W22(W22TO88), .W23(W23TO88), .W24(W24TO88), .W25(W25TO88), .W26(W26TO88), .W27(W27TO88), .W28(W28TO88), .W29(W29TO88), .W30(W30TO88), .W31(W31TO88), .W32(W32TO88), .W33(W33TO88), .W34(W34TO88), .W35(W35TO88), .W36(W36TO88), .W37(W37TO88), .W38(W38TO88), .W39(W39TO88), .W40(W40TO88), .W41(W41TO88), .W42(W42TO88), .W43(W43TO88), .W44(W44TO88), .W45(W45TO88), .W46(W46TO88), .W47(W47TO88), .W48(W48TO88), .W49(W49TO88), .W50(W50TO88), .W51(W51TO88), .W52(W52TO88), .W53(W53TO88), .W54(W54TO88), .W55(W55TO88), .W56(W56TO88), .W57(W57TO88), .W58(W58TO88), .W59(W59TO88), .W60(W60TO88), .W61(W61TO88), .W62(W62TO88), .W63(W63TO88)) neuron88(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out88));
neuron64in #(.W0(W0TO89), .W1(W1TO89), .W2(W2TO89), .W3(W3TO89), .W4(W4TO89), .W5(W5TO89), .W6(W6TO89), .W7(W7TO89), .W8(W8TO89), .W9(W9TO89), .W10(W10TO89), .W11(W11TO89), .W12(W12TO89), .W13(W13TO89), .W14(W14TO89), .W15(W15TO89), .W16(W16TO89), .W17(W17TO89), .W18(W18TO89), .W19(W19TO89), .W20(W20TO89), .W21(W21TO89), .W22(W22TO89), .W23(W23TO89), .W24(W24TO89), .W25(W25TO89), .W26(W26TO89), .W27(W27TO89), .W28(W28TO89), .W29(W29TO89), .W30(W30TO89), .W31(W31TO89), .W32(W32TO89), .W33(W33TO89), .W34(W34TO89), .W35(W35TO89), .W36(W36TO89), .W37(W37TO89), .W38(W38TO89), .W39(W39TO89), .W40(W40TO89), .W41(W41TO89), .W42(W42TO89), .W43(W43TO89), .W44(W44TO89), .W45(W45TO89), .W46(W46TO89), .W47(W47TO89), .W48(W48TO89), .W49(W49TO89), .W50(W50TO89), .W51(W51TO89), .W52(W52TO89), .W53(W53TO89), .W54(W54TO89), .W55(W55TO89), .W56(W56TO89), .W57(W57TO89), .W58(W58TO89), .W59(W59TO89), .W60(W60TO89), .W61(W61TO89), .W62(W62TO89), .W63(W63TO89)) neuron89(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out89));
neuron64in #(.W0(W0TO90), .W1(W1TO90), .W2(W2TO90), .W3(W3TO90), .W4(W4TO90), .W5(W5TO90), .W6(W6TO90), .W7(W7TO90), .W8(W8TO90), .W9(W9TO90), .W10(W10TO90), .W11(W11TO90), .W12(W12TO90), .W13(W13TO90), .W14(W14TO90), .W15(W15TO90), .W16(W16TO90), .W17(W17TO90), .W18(W18TO90), .W19(W19TO90), .W20(W20TO90), .W21(W21TO90), .W22(W22TO90), .W23(W23TO90), .W24(W24TO90), .W25(W25TO90), .W26(W26TO90), .W27(W27TO90), .W28(W28TO90), .W29(W29TO90), .W30(W30TO90), .W31(W31TO90), .W32(W32TO90), .W33(W33TO90), .W34(W34TO90), .W35(W35TO90), .W36(W36TO90), .W37(W37TO90), .W38(W38TO90), .W39(W39TO90), .W40(W40TO90), .W41(W41TO90), .W42(W42TO90), .W43(W43TO90), .W44(W44TO90), .W45(W45TO90), .W46(W46TO90), .W47(W47TO90), .W48(W48TO90), .W49(W49TO90), .W50(W50TO90), .W51(W51TO90), .W52(W52TO90), .W53(W53TO90), .W54(W54TO90), .W55(W55TO90), .W56(W56TO90), .W57(W57TO90), .W58(W58TO90), .W59(W59TO90), .W60(W60TO90), .W61(W61TO90), .W62(W62TO90), .W63(W63TO90)) neuron90(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out90));
neuron64in #(.W0(W0TO91), .W1(W1TO91), .W2(W2TO91), .W3(W3TO91), .W4(W4TO91), .W5(W5TO91), .W6(W6TO91), .W7(W7TO91), .W8(W8TO91), .W9(W9TO91), .W10(W10TO91), .W11(W11TO91), .W12(W12TO91), .W13(W13TO91), .W14(W14TO91), .W15(W15TO91), .W16(W16TO91), .W17(W17TO91), .W18(W18TO91), .W19(W19TO91), .W20(W20TO91), .W21(W21TO91), .W22(W22TO91), .W23(W23TO91), .W24(W24TO91), .W25(W25TO91), .W26(W26TO91), .W27(W27TO91), .W28(W28TO91), .W29(W29TO91), .W30(W30TO91), .W31(W31TO91), .W32(W32TO91), .W33(W33TO91), .W34(W34TO91), .W35(W35TO91), .W36(W36TO91), .W37(W37TO91), .W38(W38TO91), .W39(W39TO91), .W40(W40TO91), .W41(W41TO91), .W42(W42TO91), .W43(W43TO91), .W44(W44TO91), .W45(W45TO91), .W46(W46TO91), .W47(W47TO91), .W48(W48TO91), .W49(W49TO91), .W50(W50TO91), .W51(W51TO91), .W52(W52TO91), .W53(W53TO91), .W54(W54TO91), .W55(W55TO91), .W56(W56TO91), .W57(W57TO91), .W58(W58TO91), .W59(W59TO91), .W60(W60TO91), .W61(W61TO91), .W62(W62TO91), .W63(W63TO91)) neuron91(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out91));
neuron64in #(.W0(W0TO92), .W1(W1TO92), .W2(W2TO92), .W3(W3TO92), .W4(W4TO92), .W5(W5TO92), .W6(W6TO92), .W7(W7TO92), .W8(W8TO92), .W9(W9TO92), .W10(W10TO92), .W11(W11TO92), .W12(W12TO92), .W13(W13TO92), .W14(W14TO92), .W15(W15TO92), .W16(W16TO92), .W17(W17TO92), .W18(W18TO92), .W19(W19TO92), .W20(W20TO92), .W21(W21TO92), .W22(W22TO92), .W23(W23TO92), .W24(W24TO92), .W25(W25TO92), .W26(W26TO92), .W27(W27TO92), .W28(W28TO92), .W29(W29TO92), .W30(W30TO92), .W31(W31TO92), .W32(W32TO92), .W33(W33TO92), .W34(W34TO92), .W35(W35TO92), .W36(W36TO92), .W37(W37TO92), .W38(W38TO92), .W39(W39TO92), .W40(W40TO92), .W41(W41TO92), .W42(W42TO92), .W43(W43TO92), .W44(W44TO92), .W45(W45TO92), .W46(W46TO92), .W47(W47TO92), .W48(W48TO92), .W49(W49TO92), .W50(W50TO92), .W51(W51TO92), .W52(W52TO92), .W53(W53TO92), .W54(W54TO92), .W55(W55TO92), .W56(W56TO92), .W57(W57TO92), .W58(W58TO92), .W59(W59TO92), .W60(W60TO92), .W61(W61TO92), .W62(W62TO92), .W63(W63TO92)) neuron92(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out92));
neuron64in #(.W0(W0TO93), .W1(W1TO93), .W2(W2TO93), .W3(W3TO93), .W4(W4TO93), .W5(W5TO93), .W6(W6TO93), .W7(W7TO93), .W8(W8TO93), .W9(W9TO93), .W10(W10TO93), .W11(W11TO93), .W12(W12TO93), .W13(W13TO93), .W14(W14TO93), .W15(W15TO93), .W16(W16TO93), .W17(W17TO93), .W18(W18TO93), .W19(W19TO93), .W20(W20TO93), .W21(W21TO93), .W22(W22TO93), .W23(W23TO93), .W24(W24TO93), .W25(W25TO93), .W26(W26TO93), .W27(W27TO93), .W28(W28TO93), .W29(W29TO93), .W30(W30TO93), .W31(W31TO93), .W32(W32TO93), .W33(W33TO93), .W34(W34TO93), .W35(W35TO93), .W36(W36TO93), .W37(W37TO93), .W38(W38TO93), .W39(W39TO93), .W40(W40TO93), .W41(W41TO93), .W42(W42TO93), .W43(W43TO93), .W44(W44TO93), .W45(W45TO93), .W46(W46TO93), .W47(W47TO93), .W48(W48TO93), .W49(W49TO93), .W50(W50TO93), .W51(W51TO93), .W52(W52TO93), .W53(W53TO93), .W54(W54TO93), .W55(W55TO93), .W56(W56TO93), .W57(W57TO93), .W58(W58TO93), .W59(W59TO93), .W60(W60TO93), .W61(W61TO93), .W62(W62TO93), .W63(W63TO93)) neuron93(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out93));
neuron64in #(.W0(W0TO94), .W1(W1TO94), .W2(W2TO94), .W3(W3TO94), .W4(W4TO94), .W5(W5TO94), .W6(W6TO94), .W7(W7TO94), .W8(W8TO94), .W9(W9TO94), .W10(W10TO94), .W11(W11TO94), .W12(W12TO94), .W13(W13TO94), .W14(W14TO94), .W15(W15TO94), .W16(W16TO94), .W17(W17TO94), .W18(W18TO94), .W19(W19TO94), .W20(W20TO94), .W21(W21TO94), .W22(W22TO94), .W23(W23TO94), .W24(W24TO94), .W25(W25TO94), .W26(W26TO94), .W27(W27TO94), .W28(W28TO94), .W29(W29TO94), .W30(W30TO94), .W31(W31TO94), .W32(W32TO94), .W33(W33TO94), .W34(W34TO94), .W35(W35TO94), .W36(W36TO94), .W37(W37TO94), .W38(W38TO94), .W39(W39TO94), .W40(W40TO94), .W41(W41TO94), .W42(W42TO94), .W43(W43TO94), .W44(W44TO94), .W45(W45TO94), .W46(W46TO94), .W47(W47TO94), .W48(W48TO94), .W49(W49TO94), .W50(W50TO94), .W51(W51TO94), .W52(W52TO94), .W53(W53TO94), .W54(W54TO94), .W55(W55TO94), .W56(W56TO94), .W57(W57TO94), .W58(W58TO94), .W59(W59TO94), .W60(W60TO94), .W61(W61TO94), .W62(W62TO94), .W63(W63TO94)) neuron94(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out94));
neuron64in #(.W0(W0TO95), .W1(W1TO95), .W2(W2TO95), .W3(W3TO95), .W4(W4TO95), .W5(W5TO95), .W6(W6TO95), .W7(W7TO95), .W8(W8TO95), .W9(W9TO95), .W10(W10TO95), .W11(W11TO95), .W12(W12TO95), .W13(W13TO95), .W14(W14TO95), .W15(W15TO95), .W16(W16TO95), .W17(W17TO95), .W18(W18TO95), .W19(W19TO95), .W20(W20TO95), .W21(W21TO95), .W22(W22TO95), .W23(W23TO95), .W24(W24TO95), .W25(W25TO95), .W26(W26TO95), .W27(W27TO95), .W28(W28TO95), .W29(W29TO95), .W30(W30TO95), .W31(W31TO95), .W32(W32TO95), .W33(W33TO95), .W34(W34TO95), .W35(W35TO95), .W36(W36TO95), .W37(W37TO95), .W38(W38TO95), .W39(W39TO95), .W40(W40TO95), .W41(W41TO95), .W42(W42TO95), .W43(W43TO95), .W44(W44TO95), .W45(W45TO95), .W46(W46TO95), .W47(W47TO95), .W48(W48TO95), .W49(W49TO95), .W50(W50TO95), .W51(W51TO95), .W52(W52TO95), .W53(W53TO95), .W54(W54TO95), .W55(W55TO95), .W56(W56TO95), .W57(W57TO95), .W58(W58TO95), .W59(W59TO95), .W60(W60TO95), .W61(W61TO95), .W62(W62TO95), .W63(W63TO95)) neuron95(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out95));
neuron64in #(.W0(W0TO96), .W1(W1TO96), .W2(W2TO96), .W3(W3TO96), .W4(W4TO96), .W5(W5TO96), .W6(W6TO96), .W7(W7TO96), .W8(W8TO96), .W9(W9TO96), .W10(W10TO96), .W11(W11TO96), .W12(W12TO96), .W13(W13TO96), .W14(W14TO96), .W15(W15TO96), .W16(W16TO96), .W17(W17TO96), .W18(W18TO96), .W19(W19TO96), .W20(W20TO96), .W21(W21TO96), .W22(W22TO96), .W23(W23TO96), .W24(W24TO96), .W25(W25TO96), .W26(W26TO96), .W27(W27TO96), .W28(W28TO96), .W29(W29TO96), .W30(W30TO96), .W31(W31TO96), .W32(W32TO96), .W33(W33TO96), .W34(W34TO96), .W35(W35TO96), .W36(W36TO96), .W37(W37TO96), .W38(W38TO96), .W39(W39TO96), .W40(W40TO96), .W41(W41TO96), .W42(W42TO96), .W43(W43TO96), .W44(W44TO96), .W45(W45TO96), .W46(W46TO96), .W47(W47TO96), .W48(W48TO96), .W49(W49TO96), .W50(W50TO96), .W51(W51TO96), .W52(W52TO96), .W53(W53TO96), .W54(W54TO96), .W55(W55TO96), .W56(W56TO96), .W57(W57TO96), .W58(W58TO96), .W59(W59TO96), .W60(W60TO96), .W61(W61TO96), .W62(W62TO96), .W63(W63TO96)) neuron96(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out96));
neuron64in #(.W0(W0TO97), .W1(W1TO97), .W2(W2TO97), .W3(W3TO97), .W4(W4TO97), .W5(W5TO97), .W6(W6TO97), .W7(W7TO97), .W8(W8TO97), .W9(W9TO97), .W10(W10TO97), .W11(W11TO97), .W12(W12TO97), .W13(W13TO97), .W14(W14TO97), .W15(W15TO97), .W16(W16TO97), .W17(W17TO97), .W18(W18TO97), .W19(W19TO97), .W20(W20TO97), .W21(W21TO97), .W22(W22TO97), .W23(W23TO97), .W24(W24TO97), .W25(W25TO97), .W26(W26TO97), .W27(W27TO97), .W28(W28TO97), .W29(W29TO97), .W30(W30TO97), .W31(W31TO97), .W32(W32TO97), .W33(W33TO97), .W34(W34TO97), .W35(W35TO97), .W36(W36TO97), .W37(W37TO97), .W38(W38TO97), .W39(W39TO97), .W40(W40TO97), .W41(W41TO97), .W42(W42TO97), .W43(W43TO97), .W44(W44TO97), .W45(W45TO97), .W46(W46TO97), .W47(W47TO97), .W48(W48TO97), .W49(W49TO97), .W50(W50TO97), .W51(W51TO97), .W52(W52TO97), .W53(W53TO97), .W54(W54TO97), .W55(W55TO97), .W56(W56TO97), .W57(W57TO97), .W58(W58TO97), .W59(W59TO97), .W60(W60TO97), .W61(W61TO97), .W62(W62TO97), .W63(W63TO97)) neuron97(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out97));
neuron64in #(.W0(W0TO98), .W1(W1TO98), .W2(W2TO98), .W3(W3TO98), .W4(W4TO98), .W5(W5TO98), .W6(W6TO98), .W7(W7TO98), .W8(W8TO98), .W9(W9TO98), .W10(W10TO98), .W11(W11TO98), .W12(W12TO98), .W13(W13TO98), .W14(W14TO98), .W15(W15TO98), .W16(W16TO98), .W17(W17TO98), .W18(W18TO98), .W19(W19TO98), .W20(W20TO98), .W21(W21TO98), .W22(W22TO98), .W23(W23TO98), .W24(W24TO98), .W25(W25TO98), .W26(W26TO98), .W27(W27TO98), .W28(W28TO98), .W29(W29TO98), .W30(W30TO98), .W31(W31TO98), .W32(W32TO98), .W33(W33TO98), .W34(W34TO98), .W35(W35TO98), .W36(W36TO98), .W37(W37TO98), .W38(W38TO98), .W39(W39TO98), .W40(W40TO98), .W41(W41TO98), .W42(W42TO98), .W43(W43TO98), .W44(W44TO98), .W45(W45TO98), .W46(W46TO98), .W47(W47TO98), .W48(W48TO98), .W49(W49TO98), .W50(W50TO98), .W51(W51TO98), .W52(W52TO98), .W53(W53TO98), .W54(W54TO98), .W55(W55TO98), .W56(W56TO98), .W57(W57TO98), .W58(W58TO98), .W59(W59TO98), .W60(W60TO98), .W61(W61TO98), .W62(W62TO98), .W63(W63TO98)) neuron98(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out98));
neuron64in #(.W0(W0TO99), .W1(W1TO99), .W2(W2TO99), .W3(W3TO99), .W4(W4TO99), .W5(W5TO99), .W6(W6TO99), .W7(W7TO99), .W8(W8TO99), .W9(W9TO99), .W10(W10TO99), .W11(W11TO99), .W12(W12TO99), .W13(W13TO99), .W14(W14TO99), .W15(W15TO99), .W16(W16TO99), .W17(W17TO99), .W18(W18TO99), .W19(W19TO99), .W20(W20TO99), .W21(W21TO99), .W22(W22TO99), .W23(W23TO99), .W24(W24TO99), .W25(W25TO99), .W26(W26TO99), .W27(W27TO99), .W28(W28TO99), .W29(W29TO99), .W30(W30TO99), .W31(W31TO99), .W32(W32TO99), .W33(W33TO99), .W34(W34TO99), .W35(W35TO99), .W36(W36TO99), .W37(W37TO99), .W38(W38TO99), .W39(W39TO99), .W40(W40TO99), .W41(W41TO99), .W42(W42TO99), .W43(W43TO99), .W44(W44TO99), .W45(W45TO99), .W46(W46TO99), .W47(W47TO99), .W48(W48TO99), .W49(W49TO99), .W50(W50TO99), .W51(W51TO99), .W52(W52TO99), .W53(W53TO99), .W54(W54TO99), .W55(W55TO99), .W56(W56TO99), .W57(W57TO99), .W58(W58TO99), .W59(W59TO99), .W60(W60TO99), .W61(W61TO99), .W62(W62TO99), .W63(W63TO99)) neuron99(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out99));

endmodule

module layer100in10out(clk, rst, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85, in86, in87, in88, in89, in90, in91, in92, in93, in94, in95, in96, in97, in98, in99, out0, out1, out2, out3, out4, out5, out6, out7, out8, out9);

parameter W0TO0 = 0;
parameter W0TO1 = 0;
parameter W0TO2 = 0;
parameter W0TO3 = 0;
parameter W0TO4 = 0;
parameter W0TO5 = 0;
parameter W0TO6 = 0;
parameter W0TO7 = 0;
parameter W0TO8 = 0;
parameter W0TO9 = 0;
parameter W1TO0 = 0;
parameter W1TO1 = 0;
parameter W1TO2 = 0;
parameter W1TO3 = 0;
parameter W1TO4 = 0;
parameter W1TO5 = 0;
parameter W1TO6 = 0;
parameter W1TO7 = 0;
parameter W1TO8 = 0;
parameter W1TO9 = 0;
parameter W2TO0 = 0;
parameter W2TO1 = 0;
parameter W2TO2 = 0;
parameter W2TO3 = 0;
parameter W2TO4 = 0;
parameter W2TO5 = 0;
parameter W2TO6 = 0;
parameter W2TO7 = 0;
parameter W2TO8 = 0;
parameter W2TO9 = 0;
parameter W3TO0 = 0;
parameter W3TO1 = 0;
parameter W3TO2 = 0;
parameter W3TO3 = 0;
parameter W3TO4 = 0;
parameter W3TO5 = 0;
parameter W3TO6 = 0;
parameter W3TO7 = 0;
parameter W3TO8 = 0;
parameter W3TO9 = 0;
parameter W4TO0 = 0;
parameter W4TO1 = 0;
parameter W4TO2 = 0;
parameter W4TO3 = 0;
parameter W4TO4 = 0;
parameter W4TO5 = 0;
parameter W4TO6 = 0;
parameter W4TO7 = 0;
parameter W4TO8 = 0;
parameter W4TO9 = 0;
parameter W5TO0 = 0;
parameter W5TO1 = 0;
parameter W5TO2 = 0;
parameter W5TO3 = 0;
parameter W5TO4 = 0;
parameter W5TO5 = 0;
parameter W5TO6 = 0;
parameter W5TO7 = 0;
parameter W5TO8 = 0;
parameter W5TO9 = 0;
parameter W6TO0 = 0;
parameter W6TO1 = 0;
parameter W6TO2 = 0;
parameter W6TO3 = 0;
parameter W6TO4 = 0;
parameter W6TO5 = 0;
parameter W6TO6 = 0;
parameter W6TO7 = 0;
parameter W6TO8 = 0;
parameter W6TO9 = 0;
parameter W7TO0 = 0;
parameter W7TO1 = 0;
parameter W7TO2 = 0;
parameter W7TO3 = 0;
parameter W7TO4 = 0;
parameter W7TO5 = 0;
parameter W7TO6 = 0;
parameter W7TO7 = 0;
parameter W7TO8 = 0;
parameter W7TO9 = 0;
parameter W8TO0 = 0;
parameter W8TO1 = 0;
parameter W8TO2 = 0;
parameter W8TO3 = 0;
parameter W8TO4 = 0;
parameter W8TO5 = 0;
parameter W8TO6 = 0;
parameter W8TO7 = 0;
parameter W8TO8 = 0;
parameter W8TO9 = 0;
parameter W9TO0 = 0;
parameter W9TO1 = 0;
parameter W9TO2 = 0;
parameter W9TO3 = 0;
parameter W9TO4 = 0;
parameter W9TO5 = 0;
parameter W9TO6 = 0;
parameter W9TO7 = 0;
parameter W9TO8 = 0;
parameter W9TO9 = 0;
parameter W10TO0 = 0;
parameter W10TO1 = 0;
parameter W10TO2 = 0;
parameter W10TO3 = 0;
parameter W10TO4 = 0;
parameter W10TO5 = 0;
parameter W10TO6 = 0;
parameter W10TO7 = 0;
parameter W10TO8 = 0;
parameter W10TO9 = 0;
parameter W11TO0 = 0;
parameter W11TO1 = 0;
parameter W11TO2 = 0;
parameter W11TO3 = 0;
parameter W11TO4 = 0;
parameter W11TO5 = 0;
parameter W11TO6 = 0;
parameter W11TO7 = 0;
parameter W11TO8 = 0;
parameter W11TO9 = 0;
parameter W12TO0 = 0;
parameter W12TO1 = 0;
parameter W12TO2 = 0;
parameter W12TO3 = 0;
parameter W12TO4 = 0;
parameter W12TO5 = 0;
parameter W12TO6 = 0;
parameter W12TO7 = 0;
parameter W12TO8 = 0;
parameter W12TO9 = 0;
parameter W13TO0 = 0;
parameter W13TO1 = 0;
parameter W13TO2 = 0;
parameter W13TO3 = 0;
parameter W13TO4 = 0;
parameter W13TO5 = 0;
parameter W13TO6 = 0;
parameter W13TO7 = 0;
parameter W13TO8 = 0;
parameter W13TO9 = 0;
parameter W14TO0 = 0;
parameter W14TO1 = 0;
parameter W14TO2 = 0;
parameter W14TO3 = 0;
parameter W14TO4 = 0;
parameter W14TO5 = 0;
parameter W14TO6 = 0;
parameter W14TO7 = 0;
parameter W14TO8 = 0;
parameter W14TO9 = 0;
parameter W15TO0 = 0;
parameter W15TO1 = 0;
parameter W15TO2 = 0;
parameter W15TO3 = 0;
parameter W15TO4 = 0;
parameter W15TO5 = 0;
parameter W15TO6 = 0;
parameter W15TO7 = 0;
parameter W15TO8 = 0;
parameter W15TO9 = 0;
parameter W16TO0 = 0;
parameter W16TO1 = 0;
parameter W16TO2 = 0;
parameter W16TO3 = 0;
parameter W16TO4 = 0;
parameter W16TO5 = 0;
parameter W16TO6 = 0;
parameter W16TO7 = 0;
parameter W16TO8 = 0;
parameter W16TO9 = 0;
parameter W17TO0 = 0;
parameter W17TO1 = 0;
parameter W17TO2 = 0;
parameter W17TO3 = 0;
parameter W17TO4 = 0;
parameter W17TO5 = 0;
parameter W17TO6 = 0;
parameter W17TO7 = 0;
parameter W17TO8 = 0;
parameter W17TO9 = 0;
parameter W18TO0 = 0;
parameter W18TO1 = 0;
parameter W18TO2 = 0;
parameter W18TO3 = 0;
parameter W18TO4 = 0;
parameter W18TO5 = 0;
parameter W18TO6 = 0;
parameter W18TO7 = 0;
parameter W18TO8 = 0;
parameter W18TO9 = 0;
parameter W19TO0 = 0;
parameter W19TO1 = 0;
parameter W19TO2 = 0;
parameter W19TO3 = 0;
parameter W19TO4 = 0;
parameter W19TO5 = 0;
parameter W19TO6 = 0;
parameter W19TO7 = 0;
parameter W19TO8 = 0;
parameter W19TO9 = 0;
parameter W20TO0 = 0;
parameter W20TO1 = 0;
parameter W20TO2 = 0;
parameter W20TO3 = 0;
parameter W20TO4 = 0;
parameter W20TO5 = 0;
parameter W20TO6 = 0;
parameter W20TO7 = 0;
parameter W20TO8 = 0;
parameter W20TO9 = 0;
parameter W21TO0 = 0;
parameter W21TO1 = 0;
parameter W21TO2 = 0;
parameter W21TO3 = 0;
parameter W21TO4 = 0;
parameter W21TO5 = 0;
parameter W21TO6 = 0;
parameter W21TO7 = 0;
parameter W21TO8 = 0;
parameter W21TO9 = 0;
parameter W22TO0 = 0;
parameter W22TO1 = 0;
parameter W22TO2 = 0;
parameter W22TO3 = 0;
parameter W22TO4 = 0;
parameter W22TO5 = 0;
parameter W22TO6 = 0;
parameter W22TO7 = 0;
parameter W22TO8 = 0;
parameter W22TO9 = 0;
parameter W23TO0 = 0;
parameter W23TO1 = 0;
parameter W23TO2 = 0;
parameter W23TO3 = 0;
parameter W23TO4 = 0;
parameter W23TO5 = 0;
parameter W23TO6 = 0;
parameter W23TO7 = 0;
parameter W23TO8 = 0;
parameter W23TO9 = 0;
parameter W24TO0 = 0;
parameter W24TO1 = 0;
parameter W24TO2 = 0;
parameter W24TO3 = 0;
parameter W24TO4 = 0;
parameter W24TO5 = 0;
parameter W24TO6 = 0;
parameter W24TO7 = 0;
parameter W24TO8 = 0;
parameter W24TO9 = 0;
parameter W25TO0 = 0;
parameter W25TO1 = 0;
parameter W25TO2 = 0;
parameter W25TO3 = 0;
parameter W25TO4 = 0;
parameter W25TO5 = 0;
parameter W25TO6 = 0;
parameter W25TO7 = 0;
parameter W25TO8 = 0;
parameter W25TO9 = 0;
parameter W26TO0 = 0;
parameter W26TO1 = 0;
parameter W26TO2 = 0;
parameter W26TO3 = 0;
parameter W26TO4 = 0;
parameter W26TO5 = 0;
parameter W26TO6 = 0;
parameter W26TO7 = 0;
parameter W26TO8 = 0;
parameter W26TO9 = 0;
parameter W27TO0 = 0;
parameter W27TO1 = 0;
parameter W27TO2 = 0;
parameter W27TO3 = 0;
parameter W27TO4 = 0;
parameter W27TO5 = 0;
parameter W27TO6 = 0;
parameter W27TO7 = 0;
parameter W27TO8 = 0;
parameter W27TO9 = 0;
parameter W28TO0 = 0;
parameter W28TO1 = 0;
parameter W28TO2 = 0;
parameter W28TO3 = 0;
parameter W28TO4 = 0;
parameter W28TO5 = 0;
parameter W28TO6 = 0;
parameter W28TO7 = 0;
parameter W28TO8 = 0;
parameter W28TO9 = 0;
parameter W29TO0 = 0;
parameter W29TO1 = 0;
parameter W29TO2 = 0;
parameter W29TO3 = 0;
parameter W29TO4 = 0;
parameter W29TO5 = 0;
parameter W29TO6 = 0;
parameter W29TO7 = 0;
parameter W29TO8 = 0;
parameter W29TO9 = 0;
parameter W30TO0 = 0;
parameter W30TO1 = 0;
parameter W30TO2 = 0;
parameter W30TO3 = 0;
parameter W30TO4 = 0;
parameter W30TO5 = 0;
parameter W30TO6 = 0;
parameter W30TO7 = 0;
parameter W30TO8 = 0;
parameter W30TO9 = 0;
parameter W31TO0 = 0;
parameter W31TO1 = 0;
parameter W31TO2 = 0;
parameter W31TO3 = 0;
parameter W31TO4 = 0;
parameter W31TO5 = 0;
parameter W31TO6 = 0;
parameter W31TO7 = 0;
parameter W31TO8 = 0;
parameter W31TO9 = 0;
parameter W32TO0 = 0;
parameter W32TO1 = 0;
parameter W32TO2 = 0;
parameter W32TO3 = 0;
parameter W32TO4 = 0;
parameter W32TO5 = 0;
parameter W32TO6 = 0;
parameter W32TO7 = 0;
parameter W32TO8 = 0;
parameter W32TO9 = 0;
parameter W33TO0 = 0;
parameter W33TO1 = 0;
parameter W33TO2 = 0;
parameter W33TO3 = 0;
parameter W33TO4 = 0;
parameter W33TO5 = 0;
parameter W33TO6 = 0;
parameter W33TO7 = 0;
parameter W33TO8 = 0;
parameter W33TO9 = 0;
parameter W34TO0 = 0;
parameter W34TO1 = 0;
parameter W34TO2 = 0;
parameter W34TO3 = 0;
parameter W34TO4 = 0;
parameter W34TO5 = 0;
parameter W34TO6 = 0;
parameter W34TO7 = 0;
parameter W34TO8 = 0;
parameter W34TO9 = 0;
parameter W35TO0 = 0;
parameter W35TO1 = 0;
parameter W35TO2 = 0;
parameter W35TO3 = 0;
parameter W35TO4 = 0;
parameter W35TO5 = 0;
parameter W35TO6 = 0;
parameter W35TO7 = 0;
parameter W35TO8 = 0;
parameter W35TO9 = 0;
parameter W36TO0 = 0;
parameter W36TO1 = 0;
parameter W36TO2 = 0;
parameter W36TO3 = 0;
parameter W36TO4 = 0;
parameter W36TO5 = 0;
parameter W36TO6 = 0;
parameter W36TO7 = 0;
parameter W36TO8 = 0;
parameter W36TO9 = 0;
parameter W37TO0 = 0;
parameter W37TO1 = 0;
parameter W37TO2 = 0;
parameter W37TO3 = 0;
parameter W37TO4 = 0;
parameter W37TO5 = 0;
parameter W37TO6 = 0;
parameter W37TO7 = 0;
parameter W37TO8 = 0;
parameter W37TO9 = 0;
parameter W38TO0 = 0;
parameter W38TO1 = 0;
parameter W38TO2 = 0;
parameter W38TO3 = 0;
parameter W38TO4 = 0;
parameter W38TO5 = 0;
parameter W38TO6 = 0;
parameter W38TO7 = 0;
parameter W38TO8 = 0;
parameter W38TO9 = 0;
parameter W39TO0 = 0;
parameter W39TO1 = 0;
parameter W39TO2 = 0;
parameter W39TO3 = 0;
parameter W39TO4 = 0;
parameter W39TO5 = 0;
parameter W39TO6 = 0;
parameter W39TO7 = 0;
parameter W39TO8 = 0;
parameter W39TO9 = 0;
parameter W40TO0 = 0;
parameter W40TO1 = 0;
parameter W40TO2 = 0;
parameter W40TO3 = 0;
parameter W40TO4 = 0;
parameter W40TO5 = 0;
parameter W40TO6 = 0;
parameter W40TO7 = 0;
parameter W40TO8 = 0;
parameter W40TO9 = 0;
parameter W41TO0 = 0;
parameter W41TO1 = 0;
parameter W41TO2 = 0;
parameter W41TO3 = 0;
parameter W41TO4 = 0;
parameter W41TO5 = 0;
parameter W41TO6 = 0;
parameter W41TO7 = 0;
parameter W41TO8 = 0;
parameter W41TO9 = 0;
parameter W42TO0 = 0;
parameter W42TO1 = 0;
parameter W42TO2 = 0;
parameter W42TO3 = 0;
parameter W42TO4 = 0;
parameter W42TO5 = 0;
parameter W42TO6 = 0;
parameter W42TO7 = 0;
parameter W42TO8 = 0;
parameter W42TO9 = 0;
parameter W43TO0 = 0;
parameter W43TO1 = 0;
parameter W43TO2 = 0;
parameter W43TO3 = 0;
parameter W43TO4 = 0;
parameter W43TO5 = 0;
parameter W43TO6 = 0;
parameter W43TO7 = 0;
parameter W43TO8 = 0;
parameter W43TO9 = 0;
parameter W44TO0 = 0;
parameter W44TO1 = 0;
parameter W44TO2 = 0;
parameter W44TO3 = 0;
parameter W44TO4 = 0;
parameter W44TO5 = 0;
parameter W44TO6 = 0;
parameter W44TO7 = 0;
parameter W44TO8 = 0;
parameter W44TO9 = 0;
parameter W45TO0 = 0;
parameter W45TO1 = 0;
parameter W45TO2 = 0;
parameter W45TO3 = 0;
parameter W45TO4 = 0;
parameter W45TO5 = 0;
parameter W45TO6 = 0;
parameter W45TO7 = 0;
parameter W45TO8 = 0;
parameter W45TO9 = 0;
parameter W46TO0 = 0;
parameter W46TO1 = 0;
parameter W46TO2 = 0;
parameter W46TO3 = 0;
parameter W46TO4 = 0;
parameter W46TO5 = 0;
parameter W46TO6 = 0;
parameter W46TO7 = 0;
parameter W46TO8 = 0;
parameter W46TO9 = 0;
parameter W47TO0 = 0;
parameter W47TO1 = 0;
parameter W47TO2 = 0;
parameter W47TO3 = 0;
parameter W47TO4 = 0;
parameter W47TO5 = 0;
parameter W47TO6 = 0;
parameter W47TO7 = 0;
parameter W47TO8 = 0;
parameter W47TO9 = 0;
parameter W48TO0 = 0;
parameter W48TO1 = 0;
parameter W48TO2 = 0;
parameter W48TO3 = 0;
parameter W48TO4 = 0;
parameter W48TO5 = 0;
parameter W48TO6 = 0;
parameter W48TO7 = 0;
parameter W48TO8 = 0;
parameter W48TO9 = 0;
parameter W49TO0 = 0;
parameter W49TO1 = 0;
parameter W49TO2 = 0;
parameter W49TO3 = 0;
parameter W49TO4 = 0;
parameter W49TO5 = 0;
parameter W49TO6 = 0;
parameter W49TO7 = 0;
parameter W49TO8 = 0;
parameter W49TO9 = 0;
parameter W50TO0 = 0;
parameter W50TO1 = 0;
parameter W50TO2 = 0;
parameter W50TO3 = 0;
parameter W50TO4 = 0;
parameter W50TO5 = 0;
parameter W50TO6 = 0;
parameter W50TO7 = 0;
parameter W50TO8 = 0;
parameter W50TO9 = 0;
parameter W51TO0 = 0;
parameter W51TO1 = 0;
parameter W51TO2 = 0;
parameter W51TO3 = 0;
parameter W51TO4 = 0;
parameter W51TO5 = 0;
parameter W51TO6 = 0;
parameter W51TO7 = 0;
parameter W51TO8 = 0;
parameter W51TO9 = 0;
parameter W52TO0 = 0;
parameter W52TO1 = 0;
parameter W52TO2 = 0;
parameter W52TO3 = 0;
parameter W52TO4 = 0;
parameter W52TO5 = 0;
parameter W52TO6 = 0;
parameter W52TO7 = 0;
parameter W52TO8 = 0;
parameter W52TO9 = 0;
parameter W53TO0 = 0;
parameter W53TO1 = 0;
parameter W53TO2 = 0;
parameter W53TO3 = 0;
parameter W53TO4 = 0;
parameter W53TO5 = 0;
parameter W53TO6 = 0;
parameter W53TO7 = 0;
parameter W53TO8 = 0;
parameter W53TO9 = 0;
parameter W54TO0 = 0;
parameter W54TO1 = 0;
parameter W54TO2 = 0;
parameter W54TO3 = 0;
parameter W54TO4 = 0;
parameter W54TO5 = 0;
parameter W54TO6 = 0;
parameter W54TO7 = 0;
parameter W54TO8 = 0;
parameter W54TO9 = 0;
parameter W55TO0 = 0;
parameter W55TO1 = 0;
parameter W55TO2 = 0;
parameter W55TO3 = 0;
parameter W55TO4 = 0;
parameter W55TO5 = 0;
parameter W55TO6 = 0;
parameter W55TO7 = 0;
parameter W55TO8 = 0;
parameter W55TO9 = 0;
parameter W56TO0 = 0;
parameter W56TO1 = 0;
parameter W56TO2 = 0;
parameter W56TO3 = 0;
parameter W56TO4 = 0;
parameter W56TO5 = 0;
parameter W56TO6 = 0;
parameter W56TO7 = 0;
parameter W56TO8 = 0;
parameter W56TO9 = 0;
parameter W57TO0 = 0;
parameter W57TO1 = 0;
parameter W57TO2 = 0;
parameter W57TO3 = 0;
parameter W57TO4 = 0;
parameter W57TO5 = 0;
parameter W57TO6 = 0;
parameter W57TO7 = 0;
parameter W57TO8 = 0;
parameter W57TO9 = 0;
parameter W58TO0 = 0;
parameter W58TO1 = 0;
parameter W58TO2 = 0;
parameter W58TO3 = 0;
parameter W58TO4 = 0;
parameter W58TO5 = 0;
parameter W58TO6 = 0;
parameter W58TO7 = 0;
parameter W58TO8 = 0;
parameter W58TO9 = 0;
parameter W59TO0 = 0;
parameter W59TO1 = 0;
parameter W59TO2 = 0;
parameter W59TO3 = 0;
parameter W59TO4 = 0;
parameter W59TO5 = 0;
parameter W59TO6 = 0;
parameter W59TO7 = 0;
parameter W59TO8 = 0;
parameter W59TO9 = 0;
parameter W60TO0 = 0;
parameter W60TO1 = 0;
parameter W60TO2 = 0;
parameter W60TO3 = 0;
parameter W60TO4 = 0;
parameter W60TO5 = 0;
parameter W60TO6 = 0;
parameter W60TO7 = 0;
parameter W60TO8 = 0;
parameter W60TO9 = 0;
parameter W61TO0 = 0;
parameter W61TO1 = 0;
parameter W61TO2 = 0;
parameter W61TO3 = 0;
parameter W61TO4 = 0;
parameter W61TO5 = 0;
parameter W61TO6 = 0;
parameter W61TO7 = 0;
parameter W61TO8 = 0;
parameter W61TO9 = 0;
parameter W62TO0 = 0;
parameter W62TO1 = 0;
parameter W62TO2 = 0;
parameter W62TO3 = 0;
parameter W62TO4 = 0;
parameter W62TO5 = 0;
parameter W62TO6 = 0;
parameter W62TO7 = 0;
parameter W62TO8 = 0;
parameter W62TO9 = 0;
parameter W63TO0 = 0;
parameter W63TO1 = 0;
parameter W63TO2 = 0;
parameter W63TO3 = 0;
parameter W63TO4 = 0;
parameter W63TO5 = 0;
parameter W63TO6 = 0;
parameter W63TO7 = 0;
parameter W63TO8 = 0;
parameter W63TO9 = 0;
parameter W64TO0 = 0;
parameter W64TO1 = 0;
parameter W64TO2 = 0;
parameter W64TO3 = 0;
parameter W64TO4 = 0;
parameter W64TO5 = 0;
parameter W64TO6 = 0;
parameter W64TO7 = 0;
parameter W64TO8 = 0;
parameter W64TO9 = 0;
parameter W65TO0 = 0;
parameter W65TO1 = 0;
parameter W65TO2 = 0;
parameter W65TO3 = 0;
parameter W65TO4 = 0;
parameter W65TO5 = 0;
parameter W65TO6 = 0;
parameter W65TO7 = 0;
parameter W65TO8 = 0;
parameter W65TO9 = 0;
parameter W66TO0 = 0;
parameter W66TO1 = 0;
parameter W66TO2 = 0;
parameter W66TO3 = 0;
parameter W66TO4 = 0;
parameter W66TO5 = 0;
parameter W66TO6 = 0;
parameter W66TO7 = 0;
parameter W66TO8 = 0;
parameter W66TO9 = 0;
parameter W67TO0 = 0;
parameter W67TO1 = 0;
parameter W67TO2 = 0;
parameter W67TO3 = 0;
parameter W67TO4 = 0;
parameter W67TO5 = 0;
parameter W67TO6 = 0;
parameter W67TO7 = 0;
parameter W67TO8 = 0;
parameter W67TO9 = 0;
parameter W68TO0 = 0;
parameter W68TO1 = 0;
parameter W68TO2 = 0;
parameter W68TO3 = 0;
parameter W68TO4 = 0;
parameter W68TO5 = 0;
parameter W68TO6 = 0;
parameter W68TO7 = 0;
parameter W68TO8 = 0;
parameter W68TO9 = 0;
parameter W69TO0 = 0;
parameter W69TO1 = 0;
parameter W69TO2 = 0;
parameter W69TO3 = 0;
parameter W69TO4 = 0;
parameter W69TO5 = 0;
parameter W69TO6 = 0;
parameter W69TO7 = 0;
parameter W69TO8 = 0;
parameter W69TO9 = 0;
parameter W70TO0 = 0;
parameter W70TO1 = 0;
parameter W70TO2 = 0;
parameter W70TO3 = 0;
parameter W70TO4 = 0;
parameter W70TO5 = 0;
parameter W70TO6 = 0;
parameter W70TO7 = 0;
parameter W70TO8 = 0;
parameter W70TO9 = 0;
parameter W71TO0 = 0;
parameter W71TO1 = 0;
parameter W71TO2 = 0;
parameter W71TO3 = 0;
parameter W71TO4 = 0;
parameter W71TO5 = 0;
parameter W71TO6 = 0;
parameter W71TO7 = 0;
parameter W71TO8 = 0;
parameter W71TO9 = 0;
parameter W72TO0 = 0;
parameter W72TO1 = 0;
parameter W72TO2 = 0;
parameter W72TO3 = 0;
parameter W72TO4 = 0;
parameter W72TO5 = 0;
parameter W72TO6 = 0;
parameter W72TO7 = 0;
parameter W72TO8 = 0;
parameter W72TO9 = 0;
parameter W73TO0 = 0;
parameter W73TO1 = 0;
parameter W73TO2 = 0;
parameter W73TO3 = 0;
parameter W73TO4 = 0;
parameter W73TO5 = 0;
parameter W73TO6 = 0;
parameter W73TO7 = 0;
parameter W73TO8 = 0;
parameter W73TO9 = 0;
parameter W74TO0 = 0;
parameter W74TO1 = 0;
parameter W74TO2 = 0;
parameter W74TO3 = 0;
parameter W74TO4 = 0;
parameter W74TO5 = 0;
parameter W74TO6 = 0;
parameter W74TO7 = 0;
parameter W74TO8 = 0;
parameter W74TO9 = 0;
parameter W75TO0 = 0;
parameter W75TO1 = 0;
parameter W75TO2 = 0;
parameter W75TO3 = 0;
parameter W75TO4 = 0;
parameter W75TO5 = 0;
parameter W75TO6 = 0;
parameter W75TO7 = 0;
parameter W75TO8 = 0;
parameter W75TO9 = 0;
parameter W76TO0 = 0;
parameter W76TO1 = 0;
parameter W76TO2 = 0;
parameter W76TO3 = 0;
parameter W76TO4 = 0;
parameter W76TO5 = 0;
parameter W76TO6 = 0;
parameter W76TO7 = 0;
parameter W76TO8 = 0;
parameter W76TO9 = 0;
parameter W77TO0 = 0;
parameter W77TO1 = 0;
parameter W77TO2 = 0;
parameter W77TO3 = 0;
parameter W77TO4 = 0;
parameter W77TO5 = 0;
parameter W77TO6 = 0;
parameter W77TO7 = 0;
parameter W77TO8 = 0;
parameter W77TO9 = 0;
parameter W78TO0 = 0;
parameter W78TO1 = 0;
parameter W78TO2 = 0;
parameter W78TO3 = 0;
parameter W78TO4 = 0;
parameter W78TO5 = 0;
parameter W78TO6 = 0;
parameter W78TO7 = 0;
parameter W78TO8 = 0;
parameter W78TO9 = 0;
parameter W79TO0 = 0;
parameter W79TO1 = 0;
parameter W79TO2 = 0;
parameter W79TO3 = 0;
parameter W79TO4 = 0;
parameter W79TO5 = 0;
parameter W79TO6 = 0;
parameter W79TO7 = 0;
parameter W79TO8 = 0;
parameter W79TO9 = 0;
parameter W80TO0 = 0;
parameter W80TO1 = 0;
parameter W80TO2 = 0;
parameter W80TO3 = 0;
parameter W80TO4 = 0;
parameter W80TO5 = 0;
parameter W80TO6 = 0;
parameter W80TO7 = 0;
parameter W80TO8 = 0;
parameter W80TO9 = 0;
parameter W81TO0 = 0;
parameter W81TO1 = 0;
parameter W81TO2 = 0;
parameter W81TO3 = 0;
parameter W81TO4 = 0;
parameter W81TO5 = 0;
parameter W81TO6 = 0;
parameter W81TO7 = 0;
parameter W81TO8 = 0;
parameter W81TO9 = 0;
parameter W82TO0 = 0;
parameter W82TO1 = 0;
parameter W82TO2 = 0;
parameter W82TO3 = 0;
parameter W82TO4 = 0;
parameter W82TO5 = 0;
parameter W82TO6 = 0;
parameter W82TO7 = 0;
parameter W82TO8 = 0;
parameter W82TO9 = 0;
parameter W83TO0 = 0;
parameter W83TO1 = 0;
parameter W83TO2 = 0;
parameter W83TO3 = 0;
parameter W83TO4 = 0;
parameter W83TO5 = 0;
parameter W83TO6 = 0;
parameter W83TO7 = 0;
parameter W83TO8 = 0;
parameter W83TO9 = 0;
parameter W84TO0 = 0;
parameter W84TO1 = 0;
parameter W84TO2 = 0;
parameter W84TO3 = 0;
parameter W84TO4 = 0;
parameter W84TO5 = 0;
parameter W84TO6 = 0;
parameter W84TO7 = 0;
parameter W84TO8 = 0;
parameter W84TO9 = 0;
parameter W85TO0 = 0;
parameter W85TO1 = 0;
parameter W85TO2 = 0;
parameter W85TO3 = 0;
parameter W85TO4 = 0;
parameter W85TO5 = 0;
parameter W85TO6 = 0;
parameter W85TO7 = 0;
parameter W85TO8 = 0;
parameter W85TO9 = 0;
parameter W86TO0 = 0;
parameter W86TO1 = 0;
parameter W86TO2 = 0;
parameter W86TO3 = 0;
parameter W86TO4 = 0;
parameter W86TO5 = 0;
parameter W86TO6 = 0;
parameter W86TO7 = 0;
parameter W86TO8 = 0;
parameter W86TO9 = 0;
parameter W87TO0 = 0;
parameter W87TO1 = 0;
parameter W87TO2 = 0;
parameter W87TO3 = 0;
parameter W87TO4 = 0;
parameter W87TO5 = 0;
parameter W87TO6 = 0;
parameter W87TO7 = 0;
parameter W87TO8 = 0;
parameter W87TO9 = 0;
parameter W88TO0 = 0;
parameter W88TO1 = 0;
parameter W88TO2 = 0;
parameter W88TO3 = 0;
parameter W88TO4 = 0;
parameter W88TO5 = 0;
parameter W88TO6 = 0;
parameter W88TO7 = 0;
parameter W88TO8 = 0;
parameter W88TO9 = 0;
parameter W89TO0 = 0;
parameter W89TO1 = 0;
parameter W89TO2 = 0;
parameter W89TO3 = 0;
parameter W89TO4 = 0;
parameter W89TO5 = 0;
parameter W89TO6 = 0;
parameter W89TO7 = 0;
parameter W89TO8 = 0;
parameter W89TO9 = 0;
parameter W90TO0 = 0;
parameter W90TO1 = 0;
parameter W90TO2 = 0;
parameter W90TO3 = 0;
parameter W90TO4 = 0;
parameter W90TO5 = 0;
parameter W90TO6 = 0;
parameter W90TO7 = 0;
parameter W90TO8 = 0;
parameter W90TO9 = 0;
parameter W91TO0 = 0;
parameter W91TO1 = 0;
parameter W91TO2 = 0;
parameter W91TO3 = 0;
parameter W91TO4 = 0;
parameter W91TO5 = 0;
parameter W91TO6 = 0;
parameter W91TO7 = 0;
parameter W91TO8 = 0;
parameter W91TO9 = 0;
parameter W92TO0 = 0;
parameter W92TO1 = 0;
parameter W92TO2 = 0;
parameter W92TO3 = 0;
parameter W92TO4 = 0;
parameter W92TO5 = 0;
parameter W92TO6 = 0;
parameter W92TO7 = 0;
parameter W92TO8 = 0;
parameter W92TO9 = 0;
parameter W93TO0 = 0;
parameter W93TO1 = 0;
parameter W93TO2 = 0;
parameter W93TO3 = 0;
parameter W93TO4 = 0;
parameter W93TO5 = 0;
parameter W93TO6 = 0;
parameter W93TO7 = 0;
parameter W93TO8 = 0;
parameter W93TO9 = 0;
parameter W94TO0 = 0;
parameter W94TO1 = 0;
parameter W94TO2 = 0;
parameter W94TO3 = 0;
parameter W94TO4 = 0;
parameter W94TO5 = 0;
parameter W94TO6 = 0;
parameter W94TO7 = 0;
parameter W94TO8 = 0;
parameter W94TO9 = 0;
parameter W95TO0 = 0;
parameter W95TO1 = 0;
parameter W95TO2 = 0;
parameter W95TO3 = 0;
parameter W95TO4 = 0;
parameter W95TO5 = 0;
parameter W95TO6 = 0;
parameter W95TO7 = 0;
parameter W95TO8 = 0;
parameter W95TO9 = 0;
parameter W96TO0 = 0;
parameter W96TO1 = 0;
parameter W96TO2 = 0;
parameter W96TO3 = 0;
parameter W96TO4 = 0;
parameter W96TO5 = 0;
parameter W96TO6 = 0;
parameter W96TO7 = 0;
parameter W96TO8 = 0;
parameter W96TO9 = 0;
parameter W97TO0 = 0;
parameter W97TO1 = 0;
parameter W97TO2 = 0;
parameter W97TO3 = 0;
parameter W97TO4 = 0;
parameter W97TO5 = 0;
parameter W97TO6 = 0;
parameter W97TO7 = 0;
parameter W97TO8 = 0;
parameter W97TO9 = 0;
parameter W98TO0 = 0;
parameter W98TO1 = 0;
parameter W98TO2 = 0;
parameter W98TO3 = 0;
parameter W98TO4 = 0;
parameter W98TO5 = 0;
parameter W98TO6 = 0;
parameter W98TO7 = 0;
parameter W98TO8 = 0;
parameter W98TO9 = 0;
parameter W99TO0 = 0;
parameter W99TO1 = 0;
parameter W99TO2 = 0;
parameter W99TO3 = 0;
parameter W99TO4 = 0;
parameter W99TO5 = 0;
parameter W99TO6 = 0;
parameter W99TO7 = 0;
parameter W99TO8 = 0;
parameter W99TO9 = 0;

input wire clk;
input wire rst;

input signed [15:0] in0;
input signed [15:0] in1;
input signed [15:0] in2;
input signed [15:0] in3;
input signed [15:0] in4;
input signed [15:0] in5;
input signed [15:0] in6;
input signed [15:0] in7;
input signed [15:0] in8;
input signed [15:0] in9;
input signed [15:0] in10;
input signed [15:0] in11;
input signed [15:0] in12;
input signed [15:0] in13;
input signed [15:0] in14;
input signed [15:0] in15;
input signed [15:0] in16;
input signed [15:0] in17;
input signed [15:0] in18;
input signed [15:0] in19;
input signed [15:0] in20;
input signed [15:0] in21;
input signed [15:0] in22;
input signed [15:0] in23;
input signed [15:0] in24;
input signed [15:0] in25;
input signed [15:0] in26;
input signed [15:0] in27;
input signed [15:0] in28;
input signed [15:0] in29;
input signed [15:0] in30;
input signed [15:0] in31;
input signed [15:0] in32;
input signed [15:0] in33;
input signed [15:0] in34;
input signed [15:0] in35;
input signed [15:0] in36;
input signed [15:0] in37;
input signed [15:0] in38;
input signed [15:0] in39;
input signed [15:0] in40;
input signed [15:0] in41;
input signed [15:0] in42;
input signed [15:0] in43;
input signed [15:0] in44;
input signed [15:0] in45;
input signed [15:0] in46;
input signed [15:0] in47;
input signed [15:0] in48;
input signed [15:0] in49;
input signed [15:0] in50;
input signed [15:0] in51;
input signed [15:0] in52;
input signed [15:0] in53;
input signed [15:0] in54;
input signed [15:0] in55;
input signed [15:0] in56;
input signed [15:0] in57;
input signed [15:0] in58;
input signed [15:0] in59;
input signed [15:0] in60;
input signed [15:0] in61;
input signed [15:0] in62;
input signed [15:0] in63;
input signed [15:0] in64;
input signed [15:0] in65;
input signed [15:0] in66;
input signed [15:0] in67;
input signed [15:0] in68;
input signed [15:0] in69;
input signed [15:0] in70;
input signed [15:0] in71;
input signed [15:0] in72;
input signed [15:0] in73;
input signed [15:0] in74;
input signed [15:0] in75;
input signed [15:0] in76;
input signed [15:0] in77;
input signed [15:0] in78;
input signed [15:0] in79;
input signed [15:0] in80;
input signed [15:0] in81;
input signed [15:0] in82;
input signed [15:0] in83;
input signed [15:0] in84;
input signed [15:0] in85;
input signed [15:0] in86;
input signed [15:0] in87;
input signed [15:0] in88;
input signed [15:0] in89;
input signed [15:0] in90;
input signed [15:0] in91;
input signed [15:0] in92;
input signed [15:0] in93;
input signed [15:0] in94;
input signed [15:0] in95;
input signed [15:0] in96;
input signed [15:0] in97;
input signed [15:0] in98;
input signed [15:0] in99;

output signed [15:0] out0;
output signed [15:0] out1;
output signed [15:0] out2;
output signed [15:0] out3;
output signed [15:0] out4;
output signed [15:0] out5;
output signed [15:0] out6;
output signed [15:0] out7;
output signed [15:0] out8;
output signed [15:0] out9;

neuron100in #(.W0(W0TO0), .W1(W1TO0), .W2(W2TO0), .W3(W3TO0), .W4(W4TO0), .W5(W5TO0), .W6(W6TO0), .W7(W7TO0), .W8(W8TO0), .W9(W9TO0), .W10(W10TO0), .W11(W11TO0), .W12(W12TO0), .W13(W13TO0), .W14(W14TO0), .W15(W15TO0), .W16(W16TO0), .W17(W17TO0), .W18(W18TO0), .W19(W19TO0), .W20(W20TO0), .W21(W21TO0), .W22(W22TO0), .W23(W23TO0), .W24(W24TO0), .W25(W25TO0), .W26(W26TO0), .W27(W27TO0), .W28(W28TO0), .W29(W29TO0), .W30(W30TO0), .W31(W31TO0), .W32(W32TO0), .W33(W33TO0), .W34(W34TO0), .W35(W35TO0), .W36(W36TO0), .W37(W37TO0), .W38(W38TO0), .W39(W39TO0), .W40(W40TO0), .W41(W41TO0), .W42(W42TO0), .W43(W43TO0), .W44(W44TO0), .W45(W45TO0), .W46(W46TO0), .W47(W47TO0), .W48(W48TO0), .W49(W49TO0), .W50(W50TO0), .W51(W51TO0), .W52(W52TO0), .W53(W53TO0), .W54(W54TO0), .W55(W55TO0), .W56(W56TO0), .W57(W57TO0), .W58(W58TO0), .W59(W59TO0), .W60(W60TO0), .W61(W61TO0), .W62(W62TO0), .W63(W63TO0), .W64(W64TO0), .W65(W65TO0), .W66(W66TO0), .W67(W67TO0), .W68(W68TO0), .W69(W69TO0), .W70(W70TO0), .W71(W71TO0), .W72(W72TO0), .W73(W73TO0), .W74(W74TO0), .W75(W75TO0), .W76(W76TO0), .W77(W77TO0), .W78(W78TO0), .W79(W79TO0), .W80(W80TO0), .W81(W81TO0), .W82(W82TO0), .W83(W83TO0), .W84(W84TO0), .W85(W85TO0), .W86(W86TO0), .W87(W87TO0), .W88(W88TO0), .W89(W89TO0), .W90(W90TO0), .W91(W91TO0), .W92(W92TO0), .W93(W93TO0), .W94(W94TO0), .W95(W95TO0), .W96(W96TO0), .W97(W97TO0), .W98(W98TO0), .W99(W99TO0)) neuron0(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .in65(in65), .in66(in66), .in67(in67), .in68(in68), .in69(in69), .in70(in70), .in71(in71), .in72(in72), .in73(in73), .in74(in74), .in75(in75), .in76(in76), .in77(in77), .in78(in78), .in79(in79), .in80(in80), .in81(in81), .in82(in82), .in83(in83), .in84(in84), .in85(in85), .in86(in86), .in87(in87), .in88(in88), .in89(in89), .in90(in90), .in91(in91), .in92(in92), .in93(in93), .in94(in94), .in95(in95), .in96(in96), .in97(in97), .in98(in98), .in99(in99), .out(out0));
neuron100in #(.W0(W0TO1), .W1(W1TO1), .W2(W2TO1), .W3(W3TO1), .W4(W4TO1), .W5(W5TO1), .W6(W6TO1), .W7(W7TO1), .W8(W8TO1), .W9(W9TO1), .W10(W10TO1), .W11(W11TO1), .W12(W12TO1), .W13(W13TO1), .W14(W14TO1), .W15(W15TO1), .W16(W16TO1), .W17(W17TO1), .W18(W18TO1), .W19(W19TO1), .W20(W20TO1), .W21(W21TO1), .W22(W22TO1), .W23(W23TO1), .W24(W24TO1), .W25(W25TO1), .W26(W26TO1), .W27(W27TO1), .W28(W28TO1), .W29(W29TO1), .W30(W30TO1), .W31(W31TO1), .W32(W32TO1), .W33(W33TO1), .W34(W34TO1), .W35(W35TO1), .W36(W36TO1), .W37(W37TO1), .W38(W38TO1), .W39(W39TO1), .W40(W40TO1), .W41(W41TO1), .W42(W42TO1), .W43(W43TO1), .W44(W44TO1), .W45(W45TO1), .W46(W46TO1), .W47(W47TO1), .W48(W48TO1), .W49(W49TO1), .W50(W50TO1), .W51(W51TO1), .W52(W52TO1), .W53(W53TO1), .W54(W54TO1), .W55(W55TO1), .W56(W56TO1), .W57(W57TO1), .W58(W58TO1), .W59(W59TO1), .W60(W60TO1), .W61(W61TO1), .W62(W62TO1), .W63(W63TO1), .W64(W64TO1), .W65(W65TO1), .W66(W66TO1), .W67(W67TO1), .W68(W68TO1), .W69(W69TO1), .W70(W70TO1), .W71(W71TO1), .W72(W72TO1), .W73(W73TO1), .W74(W74TO1), .W75(W75TO1), .W76(W76TO1), .W77(W77TO1), .W78(W78TO1), .W79(W79TO1), .W80(W80TO1), .W81(W81TO1), .W82(W82TO1), .W83(W83TO1), .W84(W84TO1), .W85(W85TO1), .W86(W86TO1), .W87(W87TO1), .W88(W88TO1), .W89(W89TO1), .W90(W90TO1), .W91(W91TO1), .W92(W92TO1), .W93(W93TO1), .W94(W94TO1), .W95(W95TO1), .W96(W96TO1), .W97(W97TO1), .W98(W98TO1), .W99(W99TO1)) neuron1(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .in65(in65), .in66(in66), .in67(in67), .in68(in68), .in69(in69), .in70(in70), .in71(in71), .in72(in72), .in73(in73), .in74(in74), .in75(in75), .in76(in76), .in77(in77), .in78(in78), .in79(in79), .in80(in80), .in81(in81), .in82(in82), .in83(in83), .in84(in84), .in85(in85), .in86(in86), .in87(in87), .in88(in88), .in89(in89), .in90(in90), .in91(in91), .in92(in92), .in93(in93), .in94(in94), .in95(in95), .in96(in96), .in97(in97), .in98(in98), .in99(in99), .out(out1));
neuron100in #(.W0(W0TO2), .W1(W1TO2), .W2(W2TO2), .W3(W3TO2), .W4(W4TO2), .W5(W5TO2), .W6(W6TO2), .W7(W7TO2), .W8(W8TO2), .W9(W9TO2), .W10(W10TO2), .W11(W11TO2), .W12(W12TO2), .W13(W13TO2), .W14(W14TO2), .W15(W15TO2), .W16(W16TO2), .W17(W17TO2), .W18(W18TO2), .W19(W19TO2), .W20(W20TO2), .W21(W21TO2), .W22(W22TO2), .W23(W23TO2), .W24(W24TO2), .W25(W25TO2), .W26(W26TO2), .W27(W27TO2), .W28(W28TO2), .W29(W29TO2), .W30(W30TO2), .W31(W31TO2), .W32(W32TO2), .W33(W33TO2), .W34(W34TO2), .W35(W35TO2), .W36(W36TO2), .W37(W37TO2), .W38(W38TO2), .W39(W39TO2), .W40(W40TO2), .W41(W41TO2), .W42(W42TO2), .W43(W43TO2), .W44(W44TO2), .W45(W45TO2), .W46(W46TO2), .W47(W47TO2), .W48(W48TO2), .W49(W49TO2), .W50(W50TO2), .W51(W51TO2), .W52(W52TO2), .W53(W53TO2), .W54(W54TO2), .W55(W55TO2), .W56(W56TO2), .W57(W57TO2), .W58(W58TO2), .W59(W59TO2), .W60(W60TO2), .W61(W61TO2), .W62(W62TO2), .W63(W63TO2), .W64(W64TO2), .W65(W65TO2), .W66(W66TO2), .W67(W67TO2), .W68(W68TO2), .W69(W69TO2), .W70(W70TO2), .W71(W71TO2), .W72(W72TO2), .W73(W73TO2), .W74(W74TO2), .W75(W75TO2), .W76(W76TO2), .W77(W77TO2), .W78(W78TO2), .W79(W79TO2), .W80(W80TO2), .W81(W81TO2), .W82(W82TO2), .W83(W83TO2), .W84(W84TO2), .W85(W85TO2), .W86(W86TO2), .W87(W87TO2), .W88(W88TO2), .W89(W89TO2), .W90(W90TO2), .W91(W91TO2), .W92(W92TO2), .W93(W93TO2), .W94(W94TO2), .W95(W95TO2), .W96(W96TO2), .W97(W97TO2), .W98(W98TO2), .W99(W99TO2)) neuron2(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .in65(in65), .in66(in66), .in67(in67), .in68(in68), .in69(in69), .in70(in70), .in71(in71), .in72(in72), .in73(in73), .in74(in74), .in75(in75), .in76(in76), .in77(in77), .in78(in78), .in79(in79), .in80(in80), .in81(in81), .in82(in82), .in83(in83), .in84(in84), .in85(in85), .in86(in86), .in87(in87), .in88(in88), .in89(in89), .in90(in90), .in91(in91), .in92(in92), .in93(in93), .in94(in94), .in95(in95), .in96(in96), .in97(in97), .in98(in98), .in99(in99), .out(out2));
neuron100in #(.W0(W0TO3), .W1(W1TO3), .W2(W2TO3), .W3(W3TO3), .W4(W4TO3), .W5(W5TO3), .W6(W6TO3), .W7(W7TO3), .W8(W8TO3), .W9(W9TO3), .W10(W10TO3), .W11(W11TO3), .W12(W12TO3), .W13(W13TO3), .W14(W14TO3), .W15(W15TO3), .W16(W16TO3), .W17(W17TO3), .W18(W18TO3), .W19(W19TO3), .W20(W20TO3), .W21(W21TO3), .W22(W22TO3), .W23(W23TO3), .W24(W24TO3), .W25(W25TO3), .W26(W26TO3), .W27(W27TO3), .W28(W28TO3), .W29(W29TO3), .W30(W30TO3), .W31(W31TO3), .W32(W32TO3), .W33(W33TO3), .W34(W34TO3), .W35(W35TO3), .W36(W36TO3), .W37(W37TO3), .W38(W38TO3), .W39(W39TO3), .W40(W40TO3), .W41(W41TO3), .W42(W42TO3), .W43(W43TO3), .W44(W44TO3), .W45(W45TO3), .W46(W46TO3), .W47(W47TO3), .W48(W48TO3), .W49(W49TO3), .W50(W50TO3), .W51(W51TO3), .W52(W52TO3), .W53(W53TO3), .W54(W54TO3), .W55(W55TO3), .W56(W56TO3), .W57(W57TO3), .W58(W58TO3), .W59(W59TO3), .W60(W60TO3), .W61(W61TO3), .W62(W62TO3), .W63(W63TO3), .W64(W64TO3), .W65(W65TO3), .W66(W66TO3), .W67(W67TO3), .W68(W68TO3), .W69(W69TO3), .W70(W70TO3), .W71(W71TO3), .W72(W72TO3), .W73(W73TO3), .W74(W74TO3), .W75(W75TO3), .W76(W76TO3), .W77(W77TO3), .W78(W78TO3), .W79(W79TO3), .W80(W80TO3), .W81(W81TO3), .W82(W82TO3), .W83(W83TO3), .W84(W84TO3), .W85(W85TO3), .W86(W86TO3), .W87(W87TO3), .W88(W88TO3), .W89(W89TO3), .W90(W90TO3), .W91(W91TO3), .W92(W92TO3), .W93(W93TO3), .W94(W94TO3), .W95(W95TO3), .W96(W96TO3), .W97(W97TO3), .W98(W98TO3), .W99(W99TO3)) neuron3(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .in65(in65), .in66(in66), .in67(in67), .in68(in68), .in69(in69), .in70(in70), .in71(in71), .in72(in72), .in73(in73), .in74(in74), .in75(in75), .in76(in76), .in77(in77), .in78(in78), .in79(in79), .in80(in80), .in81(in81), .in82(in82), .in83(in83), .in84(in84), .in85(in85), .in86(in86), .in87(in87), .in88(in88), .in89(in89), .in90(in90), .in91(in91), .in92(in92), .in93(in93), .in94(in94), .in95(in95), .in96(in96), .in97(in97), .in98(in98), .in99(in99), .out(out3));
neuron100in #(.W0(W0TO4), .W1(W1TO4), .W2(W2TO4), .W3(W3TO4), .W4(W4TO4), .W5(W5TO4), .W6(W6TO4), .W7(W7TO4), .W8(W8TO4), .W9(W9TO4), .W10(W10TO4), .W11(W11TO4), .W12(W12TO4), .W13(W13TO4), .W14(W14TO4), .W15(W15TO4), .W16(W16TO4), .W17(W17TO4), .W18(W18TO4), .W19(W19TO4), .W20(W20TO4), .W21(W21TO4), .W22(W22TO4), .W23(W23TO4), .W24(W24TO4), .W25(W25TO4), .W26(W26TO4), .W27(W27TO4), .W28(W28TO4), .W29(W29TO4), .W30(W30TO4), .W31(W31TO4), .W32(W32TO4), .W33(W33TO4), .W34(W34TO4), .W35(W35TO4), .W36(W36TO4), .W37(W37TO4), .W38(W38TO4), .W39(W39TO4), .W40(W40TO4), .W41(W41TO4), .W42(W42TO4), .W43(W43TO4), .W44(W44TO4), .W45(W45TO4), .W46(W46TO4), .W47(W47TO4), .W48(W48TO4), .W49(W49TO4), .W50(W50TO4), .W51(W51TO4), .W52(W52TO4), .W53(W53TO4), .W54(W54TO4), .W55(W55TO4), .W56(W56TO4), .W57(W57TO4), .W58(W58TO4), .W59(W59TO4), .W60(W60TO4), .W61(W61TO4), .W62(W62TO4), .W63(W63TO4), .W64(W64TO4), .W65(W65TO4), .W66(W66TO4), .W67(W67TO4), .W68(W68TO4), .W69(W69TO4), .W70(W70TO4), .W71(W71TO4), .W72(W72TO4), .W73(W73TO4), .W74(W74TO4), .W75(W75TO4), .W76(W76TO4), .W77(W77TO4), .W78(W78TO4), .W79(W79TO4), .W80(W80TO4), .W81(W81TO4), .W82(W82TO4), .W83(W83TO4), .W84(W84TO4), .W85(W85TO4), .W86(W86TO4), .W87(W87TO4), .W88(W88TO4), .W89(W89TO4), .W90(W90TO4), .W91(W91TO4), .W92(W92TO4), .W93(W93TO4), .W94(W94TO4), .W95(W95TO4), .W96(W96TO4), .W97(W97TO4), .W98(W98TO4), .W99(W99TO4)) neuron4(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .in65(in65), .in66(in66), .in67(in67), .in68(in68), .in69(in69), .in70(in70), .in71(in71), .in72(in72), .in73(in73), .in74(in74), .in75(in75), .in76(in76), .in77(in77), .in78(in78), .in79(in79), .in80(in80), .in81(in81), .in82(in82), .in83(in83), .in84(in84), .in85(in85), .in86(in86), .in87(in87), .in88(in88), .in89(in89), .in90(in90), .in91(in91), .in92(in92), .in93(in93), .in94(in94), .in95(in95), .in96(in96), .in97(in97), .in98(in98), .in99(in99), .out(out4));
neuron100in #(.W0(W0TO5), .W1(W1TO5), .W2(W2TO5), .W3(W3TO5), .W4(W4TO5), .W5(W5TO5), .W6(W6TO5), .W7(W7TO5), .W8(W8TO5), .W9(W9TO5), .W10(W10TO5), .W11(W11TO5), .W12(W12TO5), .W13(W13TO5), .W14(W14TO5), .W15(W15TO5), .W16(W16TO5), .W17(W17TO5), .W18(W18TO5), .W19(W19TO5), .W20(W20TO5), .W21(W21TO5), .W22(W22TO5), .W23(W23TO5), .W24(W24TO5), .W25(W25TO5), .W26(W26TO5), .W27(W27TO5), .W28(W28TO5), .W29(W29TO5), .W30(W30TO5), .W31(W31TO5), .W32(W32TO5), .W33(W33TO5), .W34(W34TO5), .W35(W35TO5), .W36(W36TO5), .W37(W37TO5), .W38(W38TO5), .W39(W39TO5), .W40(W40TO5), .W41(W41TO5), .W42(W42TO5), .W43(W43TO5), .W44(W44TO5), .W45(W45TO5), .W46(W46TO5), .W47(W47TO5), .W48(W48TO5), .W49(W49TO5), .W50(W50TO5), .W51(W51TO5), .W52(W52TO5), .W53(W53TO5), .W54(W54TO5), .W55(W55TO5), .W56(W56TO5), .W57(W57TO5), .W58(W58TO5), .W59(W59TO5), .W60(W60TO5), .W61(W61TO5), .W62(W62TO5), .W63(W63TO5), .W64(W64TO5), .W65(W65TO5), .W66(W66TO5), .W67(W67TO5), .W68(W68TO5), .W69(W69TO5), .W70(W70TO5), .W71(W71TO5), .W72(W72TO5), .W73(W73TO5), .W74(W74TO5), .W75(W75TO5), .W76(W76TO5), .W77(W77TO5), .W78(W78TO5), .W79(W79TO5), .W80(W80TO5), .W81(W81TO5), .W82(W82TO5), .W83(W83TO5), .W84(W84TO5), .W85(W85TO5), .W86(W86TO5), .W87(W87TO5), .W88(W88TO5), .W89(W89TO5), .W90(W90TO5), .W91(W91TO5), .W92(W92TO5), .W93(W93TO5), .W94(W94TO5), .W95(W95TO5), .W96(W96TO5), .W97(W97TO5), .W98(W98TO5), .W99(W99TO5)) neuron5(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .in65(in65), .in66(in66), .in67(in67), .in68(in68), .in69(in69), .in70(in70), .in71(in71), .in72(in72), .in73(in73), .in74(in74), .in75(in75), .in76(in76), .in77(in77), .in78(in78), .in79(in79), .in80(in80), .in81(in81), .in82(in82), .in83(in83), .in84(in84), .in85(in85), .in86(in86), .in87(in87), .in88(in88), .in89(in89), .in90(in90), .in91(in91), .in92(in92), .in93(in93), .in94(in94), .in95(in95), .in96(in96), .in97(in97), .in98(in98), .in99(in99), .out(out5));
neuron100in #(.W0(W0TO6), .W1(W1TO6), .W2(W2TO6), .W3(W3TO6), .W4(W4TO6), .W5(W5TO6), .W6(W6TO6), .W7(W7TO6), .W8(W8TO6), .W9(W9TO6), .W10(W10TO6), .W11(W11TO6), .W12(W12TO6), .W13(W13TO6), .W14(W14TO6), .W15(W15TO6), .W16(W16TO6), .W17(W17TO6), .W18(W18TO6), .W19(W19TO6), .W20(W20TO6), .W21(W21TO6), .W22(W22TO6), .W23(W23TO6), .W24(W24TO6), .W25(W25TO6), .W26(W26TO6), .W27(W27TO6), .W28(W28TO6), .W29(W29TO6), .W30(W30TO6), .W31(W31TO6), .W32(W32TO6), .W33(W33TO6), .W34(W34TO6), .W35(W35TO6), .W36(W36TO6), .W37(W37TO6), .W38(W38TO6), .W39(W39TO6), .W40(W40TO6), .W41(W41TO6), .W42(W42TO6), .W43(W43TO6), .W44(W44TO6), .W45(W45TO6), .W46(W46TO6), .W47(W47TO6), .W48(W48TO6), .W49(W49TO6), .W50(W50TO6), .W51(W51TO6), .W52(W52TO6), .W53(W53TO6), .W54(W54TO6), .W55(W55TO6), .W56(W56TO6), .W57(W57TO6), .W58(W58TO6), .W59(W59TO6), .W60(W60TO6), .W61(W61TO6), .W62(W62TO6), .W63(W63TO6), .W64(W64TO6), .W65(W65TO6), .W66(W66TO6), .W67(W67TO6), .W68(W68TO6), .W69(W69TO6), .W70(W70TO6), .W71(W71TO6), .W72(W72TO6), .W73(W73TO6), .W74(W74TO6), .W75(W75TO6), .W76(W76TO6), .W77(W77TO6), .W78(W78TO6), .W79(W79TO6), .W80(W80TO6), .W81(W81TO6), .W82(W82TO6), .W83(W83TO6), .W84(W84TO6), .W85(W85TO6), .W86(W86TO6), .W87(W87TO6), .W88(W88TO6), .W89(W89TO6), .W90(W90TO6), .W91(W91TO6), .W92(W92TO6), .W93(W93TO6), .W94(W94TO6), .W95(W95TO6), .W96(W96TO6), .W97(W97TO6), .W98(W98TO6), .W99(W99TO6)) neuron6(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .in65(in65), .in66(in66), .in67(in67), .in68(in68), .in69(in69), .in70(in70), .in71(in71), .in72(in72), .in73(in73), .in74(in74), .in75(in75), .in76(in76), .in77(in77), .in78(in78), .in79(in79), .in80(in80), .in81(in81), .in82(in82), .in83(in83), .in84(in84), .in85(in85), .in86(in86), .in87(in87), .in88(in88), .in89(in89), .in90(in90), .in91(in91), .in92(in92), .in93(in93), .in94(in94), .in95(in95), .in96(in96), .in97(in97), .in98(in98), .in99(in99), .out(out6));
neuron100in #(.W0(W0TO7), .W1(W1TO7), .W2(W2TO7), .W3(W3TO7), .W4(W4TO7), .W5(W5TO7), .W6(W6TO7), .W7(W7TO7), .W8(W8TO7), .W9(W9TO7), .W10(W10TO7), .W11(W11TO7), .W12(W12TO7), .W13(W13TO7), .W14(W14TO7), .W15(W15TO7), .W16(W16TO7), .W17(W17TO7), .W18(W18TO7), .W19(W19TO7), .W20(W20TO7), .W21(W21TO7), .W22(W22TO7), .W23(W23TO7), .W24(W24TO7), .W25(W25TO7), .W26(W26TO7), .W27(W27TO7), .W28(W28TO7), .W29(W29TO7), .W30(W30TO7), .W31(W31TO7), .W32(W32TO7), .W33(W33TO7), .W34(W34TO7), .W35(W35TO7), .W36(W36TO7), .W37(W37TO7), .W38(W38TO7), .W39(W39TO7), .W40(W40TO7), .W41(W41TO7), .W42(W42TO7), .W43(W43TO7), .W44(W44TO7), .W45(W45TO7), .W46(W46TO7), .W47(W47TO7), .W48(W48TO7), .W49(W49TO7), .W50(W50TO7), .W51(W51TO7), .W52(W52TO7), .W53(W53TO7), .W54(W54TO7), .W55(W55TO7), .W56(W56TO7), .W57(W57TO7), .W58(W58TO7), .W59(W59TO7), .W60(W60TO7), .W61(W61TO7), .W62(W62TO7), .W63(W63TO7), .W64(W64TO7), .W65(W65TO7), .W66(W66TO7), .W67(W67TO7), .W68(W68TO7), .W69(W69TO7), .W70(W70TO7), .W71(W71TO7), .W72(W72TO7), .W73(W73TO7), .W74(W74TO7), .W75(W75TO7), .W76(W76TO7), .W77(W77TO7), .W78(W78TO7), .W79(W79TO7), .W80(W80TO7), .W81(W81TO7), .W82(W82TO7), .W83(W83TO7), .W84(W84TO7), .W85(W85TO7), .W86(W86TO7), .W87(W87TO7), .W88(W88TO7), .W89(W89TO7), .W90(W90TO7), .W91(W91TO7), .W92(W92TO7), .W93(W93TO7), .W94(W94TO7), .W95(W95TO7), .W96(W96TO7), .W97(W97TO7), .W98(W98TO7), .W99(W99TO7)) neuron7(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .in65(in65), .in66(in66), .in67(in67), .in68(in68), .in69(in69), .in70(in70), .in71(in71), .in72(in72), .in73(in73), .in74(in74), .in75(in75), .in76(in76), .in77(in77), .in78(in78), .in79(in79), .in80(in80), .in81(in81), .in82(in82), .in83(in83), .in84(in84), .in85(in85), .in86(in86), .in87(in87), .in88(in88), .in89(in89), .in90(in90), .in91(in91), .in92(in92), .in93(in93), .in94(in94), .in95(in95), .in96(in96), .in97(in97), .in98(in98), .in99(in99), .out(out7));
neuron100in #(.W0(W0TO8), .W1(W1TO8), .W2(W2TO8), .W3(W3TO8), .W4(W4TO8), .W5(W5TO8), .W6(W6TO8), .W7(W7TO8), .W8(W8TO8), .W9(W9TO8), .W10(W10TO8), .W11(W11TO8), .W12(W12TO8), .W13(W13TO8), .W14(W14TO8), .W15(W15TO8), .W16(W16TO8), .W17(W17TO8), .W18(W18TO8), .W19(W19TO8), .W20(W20TO8), .W21(W21TO8), .W22(W22TO8), .W23(W23TO8), .W24(W24TO8), .W25(W25TO8), .W26(W26TO8), .W27(W27TO8), .W28(W28TO8), .W29(W29TO8), .W30(W30TO8), .W31(W31TO8), .W32(W32TO8), .W33(W33TO8), .W34(W34TO8), .W35(W35TO8), .W36(W36TO8), .W37(W37TO8), .W38(W38TO8), .W39(W39TO8), .W40(W40TO8), .W41(W41TO8), .W42(W42TO8), .W43(W43TO8), .W44(W44TO8), .W45(W45TO8), .W46(W46TO8), .W47(W47TO8), .W48(W48TO8), .W49(W49TO8), .W50(W50TO8), .W51(W51TO8), .W52(W52TO8), .W53(W53TO8), .W54(W54TO8), .W55(W55TO8), .W56(W56TO8), .W57(W57TO8), .W58(W58TO8), .W59(W59TO8), .W60(W60TO8), .W61(W61TO8), .W62(W62TO8), .W63(W63TO8), .W64(W64TO8), .W65(W65TO8), .W66(W66TO8), .W67(W67TO8), .W68(W68TO8), .W69(W69TO8), .W70(W70TO8), .W71(W71TO8), .W72(W72TO8), .W73(W73TO8), .W74(W74TO8), .W75(W75TO8), .W76(W76TO8), .W77(W77TO8), .W78(W78TO8), .W79(W79TO8), .W80(W80TO8), .W81(W81TO8), .W82(W82TO8), .W83(W83TO8), .W84(W84TO8), .W85(W85TO8), .W86(W86TO8), .W87(W87TO8), .W88(W88TO8), .W89(W89TO8), .W90(W90TO8), .W91(W91TO8), .W92(W92TO8), .W93(W93TO8), .W94(W94TO8), .W95(W95TO8), .W96(W96TO8), .W97(W97TO8), .W98(W98TO8), .W99(W99TO8)) neuron8(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .in65(in65), .in66(in66), .in67(in67), .in68(in68), .in69(in69), .in70(in70), .in71(in71), .in72(in72), .in73(in73), .in74(in74), .in75(in75), .in76(in76), .in77(in77), .in78(in78), .in79(in79), .in80(in80), .in81(in81), .in82(in82), .in83(in83), .in84(in84), .in85(in85), .in86(in86), .in87(in87), .in88(in88), .in89(in89), .in90(in90), .in91(in91), .in92(in92), .in93(in93), .in94(in94), .in95(in95), .in96(in96), .in97(in97), .in98(in98), .in99(in99), .out(out8));
neuron100in #(.W0(W0TO9), .W1(W1TO9), .W2(W2TO9), .W3(W3TO9), .W4(W4TO9), .W5(W5TO9), .W6(W6TO9), .W7(W7TO9), .W8(W8TO9), .W9(W9TO9), .W10(W10TO9), .W11(W11TO9), .W12(W12TO9), .W13(W13TO9), .W14(W14TO9), .W15(W15TO9), .W16(W16TO9), .W17(W17TO9), .W18(W18TO9), .W19(W19TO9), .W20(W20TO9), .W21(W21TO9), .W22(W22TO9), .W23(W23TO9), .W24(W24TO9), .W25(W25TO9), .W26(W26TO9), .W27(W27TO9), .W28(W28TO9), .W29(W29TO9), .W30(W30TO9), .W31(W31TO9), .W32(W32TO9), .W33(W33TO9), .W34(W34TO9), .W35(W35TO9), .W36(W36TO9), .W37(W37TO9), .W38(W38TO9), .W39(W39TO9), .W40(W40TO9), .W41(W41TO9), .W42(W42TO9), .W43(W43TO9), .W44(W44TO9), .W45(W45TO9), .W46(W46TO9), .W47(W47TO9), .W48(W48TO9), .W49(W49TO9), .W50(W50TO9), .W51(W51TO9), .W52(W52TO9), .W53(W53TO9), .W54(W54TO9), .W55(W55TO9), .W56(W56TO9), .W57(W57TO9), .W58(W58TO9), .W59(W59TO9), .W60(W60TO9), .W61(W61TO9), .W62(W62TO9), .W63(W63TO9), .W64(W64TO9), .W65(W65TO9), .W66(W66TO9), .W67(W67TO9), .W68(W68TO9), .W69(W69TO9), .W70(W70TO9), .W71(W71TO9), .W72(W72TO9), .W73(W73TO9), .W74(W74TO9), .W75(W75TO9), .W76(W76TO9), .W77(W77TO9), .W78(W78TO9), .W79(W79TO9), .W80(W80TO9), .W81(W81TO9), .W82(W82TO9), .W83(W83TO9), .W84(W84TO9), .W85(W85TO9), .W86(W86TO9), .W87(W87TO9), .W88(W88TO9), .W89(W89TO9), .W90(W90TO9), .W91(W91TO9), .W92(W92TO9), .W93(W93TO9), .W94(W94TO9), .W95(W95TO9), .W96(W96TO9), .W97(W97TO9), .W98(W98TO9), .W99(W99TO9)) neuron9(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .in65(in65), .in66(in66), .in67(in67), .in68(in68), .in69(in69), .in70(in70), .in71(in71), .in72(in72), .in73(in73), .in74(in74), .in75(in75), .in76(in76), .in77(in77), .in78(in78), .in79(in79), .in80(in80), .in81(in81), .in82(in82), .in83(in83), .in84(in84), .in85(in85), .in86(in86), .in87(in87), .in88(in88), .in89(in89), .in90(in90), .in91(in91), .in92(in92), .in93(in93), .in94(in94), .in95(in95), .in96(in96), .in97(in97), .in98(in98), .in99(in99), .out(out9));

endmodule

module network(clk, rst, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, out0, out1, out2, out3, out4, out5, out6, out7, out8, out9);

input wire clk;
input wire rst;

input signed [15:0] in0;
input signed [15:0] in1;
input signed [15:0] in2;
input signed [15:0] in3;
input signed [15:0] in4;
input signed [15:0] in5;
input signed [15:0] in6;
input signed [15:0] in7;
input signed [15:0] in8;
input signed [15:0] in9;
input signed [15:0] in10;
input signed [15:0] in11;
input signed [15:0] in12;
input signed [15:0] in13;
input signed [15:0] in14;
input signed [15:0] in15;
input signed [15:0] in16;
input signed [15:0] in17;
input signed [15:0] in18;
input signed [15:0] in19;
input signed [15:0] in20;
input signed [15:0] in21;
input signed [15:0] in22;
input signed [15:0] in23;
input signed [15:0] in24;
input signed [15:0] in25;
input signed [15:0] in26;
input signed [15:0] in27;
input signed [15:0] in28;
input signed [15:0] in29;
input signed [15:0] in30;
input signed [15:0] in31;
input signed [15:0] in32;
input signed [15:0] in33;
input signed [15:0] in34;
input signed [15:0] in35;
input signed [15:0] in36;
input signed [15:0] in37;
input signed [15:0] in38;
input signed [15:0] in39;
input signed [15:0] in40;
input signed [15:0] in41;
input signed [15:0] in42;
input signed [15:0] in43;
input signed [15:0] in44;
input signed [15:0] in45;
input signed [15:0] in46;
input signed [15:0] in47;
input signed [15:0] in48;
input signed [15:0] in49;
input signed [15:0] in50;
input signed [15:0] in51;
input signed [15:0] in52;
input signed [15:0] in53;
input signed [15:0] in54;
input signed [15:0] in55;
input signed [15:0] in56;
input signed [15:0] in57;
input signed [15:0] in58;
input signed [15:0] in59;
input signed [15:0] in60;
input signed [15:0] in61;
input signed [15:0] in62;
input signed [15:0] in63;

output signed [15:0] out0;
output signed [15:0] out1;
output signed [15:0] out2;
output signed [15:0] out3;
output signed [15:0] out4;
output signed [15:0] out5;
output signed [15:0] out6;
output signed [15:0] out7;
output signed [15:0] out8;
output signed [15:0] out9;

wire[15:0] con0[0:99];

layer64in100out #(.W0TO0(-14558), .W0TO1(7573), .W0TO2(11443), .W0TO3(-2290), .W0TO4(-12746), .W0TO5(8610), .W0TO6(-15647), .W0TO7(14623), .W0TO8(18759), .W0TO9(-3193), .W0TO10(5357), .W0TO11(7244), .W0TO12(-12547), .W0TO13(-18787), .W0TO14(-15874), .W0TO15(-1513), .W0TO16(16707), .W0TO17(4008), .W0TO18(-16687), .W0TO19(-17181), .W0TO20(6662), .W0TO21(-18343), .W0TO22(4320), .W0TO23(-8484), .W0TO24(10203), .W0TO25(482), .W0TO26(2474), .W0TO27(-17088), .W0TO28(8299), .W0TO29(847), .W0TO30(-9527), .W0TO31(-15259), .W0TO32(-4577), .W0TO33(-17706), .W0TO34(3095), .W0TO35(9508), .W0TO36(294), .W0TO37(-16578), .W0TO38(-17979), .W0TO39(4797), .W0TO40(11674), .W0TO41(-15791), .W0TO42(2063), .W0TO43(3410), .W0TO44(-1797), .W0TO45(2333), .W0TO46(-7386), .W0TO47(659), .W0TO48(-8241), .W0TO49(14057), .W0TO50(-14676), .W0TO51(-14885), .W0TO52(-11396), .W0TO53(10789), .W0TO54(2954), .W0TO55(11786), .W0TO56(7488), .W0TO57(10064), .W0TO58(8663), .W0TO59(6332), .W0TO60(-18780), .W0TO61(3080), .W0TO62(-4728), .W0TO63(8170), .W0TO64(3335), .W0TO65(2638), .W0TO66(9045), .W0TO67(179), .W0TO68(12021), .W0TO69(2877), .W0TO70(-16400), .W0TO71(13801), .W0TO72(-18957), .W0TO73(-8611), .W0TO74(-10688), .W0TO75(17351), .W0TO76(8167), .W0TO77(-5303), .W0TO78(3480), .W0TO79(10063), .W0TO80(-9155), .W0TO81(1668), .W0TO82(-404), .W0TO83(-1113), .W0TO84(-9920), .W0TO85(2017), .W0TO86(-11217), .W0TO87(-4284), .W0TO88(8507), .W0TO89(9673), .W0TO90(5756), .W0TO91(-6280), .W0TO92(-10310), .W0TO93(-18280), .W0TO94(11313), .W0TO95(11827), .W0TO96(11887), .W0TO97(-14042), .W0TO98(-8825), .W0TO99(-5702), .W1TO0(-15502), .W1TO1(17717), .W1TO2(8708), .W1TO3(-16448), .W1TO4(-18796), .W1TO5(-17259), .W1TO6(-1870), .W1TO7(-15047), .W1TO8(13558), .W1TO9(-15177), .W1TO10(9043), .W1TO11(-17131), .W1TO12(14930), .W1TO13(-10317), .W1TO14(-5704), .W1TO15(1326), .W1TO16(-4192), .W1TO17(-15379), .W1TO18(-6940), .W1TO19(8662), .W1TO20(-9679), .W1TO21(16226), .W1TO22(18068), .W1TO23(-18183), .W1TO24(2937), .W1TO25(-12439), .W1TO26(3593), .W1TO27(13008), .W1TO28(5693), .W1TO29(5225), .W1TO30(914), .W1TO31(-1638), .W1TO32(-9330), .W1TO33(9835), .W1TO34(9921), .W1TO35(10253), .W1TO36(-19814), .W1TO37(1831), .W1TO38(-9762), .W1TO39(-12783), .W1TO40(-11109), .W1TO41(-1203), .W1TO42(-17356), .W1TO43(-1384), .W1TO44(-13614), .W1TO45(-15432), .W1TO46(-8124), .W1TO47(-11675), .W1TO48(6369), .W1TO49(11798), .W1TO50(-10062), .W1TO51(-8057), .W1TO52(-12749), .W1TO53(16158), .W1TO54(-10175), .W1TO55(12627), .W1TO56(7029), .W1TO57(18187), .W1TO58(-14597), .W1TO59(2246), .W1TO60(7627), .W1TO61(13723), .W1TO62(14375), .W1TO63(10571), .W1TO64(5829), .W1TO65(4109), .W1TO66(7363), .W1TO67(-11880), .W1TO68(-12405), .W1TO69(10), .W1TO70(18539), .W1TO71(-2831), .W1TO72(10030), .W1TO73(-8345), .W1TO74(-18414), .W1TO75(18154), .W1TO76(6941), .W1TO77(4499), .W1TO78(15785), .W1TO79(13304), .W1TO80(-14361), .W1TO81(-15579), .W1TO82(-84), .W1TO83(18978), .W1TO84(2650), .W1TO85(2584), .W1TO86(15691), .W1TO87(-5126), .W1TO88(-10080), .W1TO89(18618), .W1TO90(13361), .W1TO91(-538), .W1TO92(-10424), .W1TO93(-8008), .W1TO94(14840), .W1TO95(7466), .W1TO96(-17947), .W1TO97(-3892), .W1TO98(-1396), .W1TO99(-11251), .W2TO0(11094), .W2TO1(7977), .W2TO2(-6201), .W2TO3(-7796), .W2TO4(8999), .W2TO5(12665), .W2TO6(17113), .W2TO7(831), .W2TO8(-12694), .W2TO9(12436), .W2TO10(-16511), .W2TO11(13200), .W2TO12(20441), .W2TO13(18039), .W2TO14(17483), .W2TO15(-15309), .W2TO16(-8458), .W2TO17(-12901), .W2TO18(-11660), .W2TO19(-4064), .W2TO20(10428), .W2TO21(7373), .W2TO22(-9797), .W2TO23(-3900), .W2TO24(-357), .W2TO25(-16336), .W2TO26(297), .W2TO27(12308), .W2TO28(78), .W2TO29(-1483), .W2TO30(-18880), .W2TO31(-48), .W2TO32(-3200), .W2TO33(10195), .W2TO34(-17669), .W2TO35(12543), .W2TO36(1550), .W2TO37(423), .W2TO38(12738), .W2TO39(3660), .W2TO40(-12810), .W2TO41(11056), .W2TO42(8259), .W2TO43(-2072), .W2TO44(-2764), .W2TO45(9017), .W2TO46(13914), .W2TO47(-15750), .W2TO48(2964), .W2TO49(-3412), .W2TO50(-8023), .W2TO51(-610), .W2TO52(18355), .W2TO53(16888), .W2TO54(4724), .W2TO55(1379), .W2TO56(1162), .W2TO57(-13965), .W2TO58(13149), .W2TO59(-7497), .W2TO60(-9932), .W2TO61(-4306), .W2TO62(-5117), .W2TO63(13797), .W2TO64(5855), .W2TO65(300), .W2TO66(14196), .W2TO67(-2025), .W2TO68(12596), .W2TO69(2882), .W2TO70(-17750), .W2TO71(10525), .W2TO72(-16822), .W2TO73(4905), .W2TO74(-8788), .W2TO75(-9610), .W2TO76(2839), .W2TO77(-9468), .W2TO78(-4739), .W2TO79(-14527), .W2TO80(4317), .W2TO81(2976), .W2TO82(-81), .W2TO83(-2602), .W2TO84(-7867), .W2TO85(6147), .W2TO86(13955), .W2TO87(557), .W2TO88(-24504), .W2TO89(-6792), .W2TO90(1416), .W2TO91(-8408), .W2TO92(-9766), .W2TO93(-7790), .W2TO94(7753), .W2TO95(3816), .W2TO96(19441), .W2TO97(14505), .W2TO98(-16336), .W2TO99(-9528), .W3TO0(-9919), .W3TO1(-17796), .W3TO2(-17121), .W3TO3(-5701), .W3TO4(17075), .W3TO5(-16561), .W3TO6(11270), .W3TO7(17902), .W3TO8(-8537), .W3TO9(12172), .W3TO10(-8812), .W3TO11(-9461), .W3TO12(-8149), .W3TO13(9578), .W3TO14(-17162), .W3TO15(-14470), .W3TO16(-12364), .W3TO17(9722), .W3TO18(1138), .W3TO19(-18135), .W3TO20(-9641), .W3TO21(-11517), .W3TO22(-14769), .W3TO23(-21238), .W3TO24(-11257), .W3TO25(-9107), .W3TO26(-12179), .W3TO27(-3205), .W3TO28(-3700), .W3TO29(218), .W3TO30(-14922), .W3TO31(-7627), .W3TO32(15609), .W3TO33(-9374), .W3TO34(7281), .W3TO35(10598), .W3TO36(12138), .W3TO37(-2093), .W3TO38(3707), .W3TO39(-20650), .W3TO40(-22029), .W3TO41(-19803), .W3TO42(-16582), .W3TO43(26), .W3TO44(-12734), .W3TO45(-11256), .W3TO46(-6009), .W3TO47(1172), .W3TO48(-1752), .W3TO49(4486), .W3TO50(17359), .W3TO51(-11056), .W3TO52(-13764), .W3TO53(12870), .W3TO54(-4860), .W3TO55(-20089), .W3TO56(-1037), .W3TO57(5855), .W3TO58(6067), .W3TO59(15317), .W3TO60(-21512), .W3TO61(2920), .W3TO62(-881), .W3TO63(21671), .W3TO64(-9045), .W3TO65(-14404), .W3TO66(5343), .W3TO67(-8041), .W3TO68(9164), .W3TO69(1314), .W3TO70(-10631), .W3TO71(15100), .W3TO72(-348), .W3TO73(-754), .W3TO74(-12741), .W3TO75(14355), .W3TO76(13225), .W3TO77(-4678), .W3TO78(4933), .W3TO79(15413), .W3TO80(-19809), .W3TO81(16809), .W3TO82(-10200), .W3TO83(11649), .W3TO84(13279), .W3TO85(18105), .W3TO86(12224), .W3TO87(-19632), .W3TO88(-4125), .W3TO89(19711), .W3TO90(11828), .W3TO91(-13822), .W3TO92(-14344), .W3TO93(-10764), .W3TO94(-2937), .W3TO95(1228), .W3TO96(13801), .W3TO97(4603), .W3TO98(12855), .W3TO99(9259), .W4TO0(13710), .W4TO1(19724), .W4TO2(6605), .W4TO3(15149), .W4TO4(-4098), .W4TO5(1603), .W4TO6(20276), .W4TO7(-3132), .W4TO8(8675), .W4TO9(-8600), .W4TO10(-6518), .W4TO11(5972), .W4TO12(4625), .W4TO13(-5355), .W4TO14(17101), .W4TO15(-10659), .W4TO16(-14858), .W4TO17(-4063), .W4TO18(12720), .W4TO19(-3772), .W4TO20(-14286), .W4TO21(-15421), .W4TO22(10306), .W4TO23(-431), .W4TO24(7054), .W4TO25(10827), .W4TO26(1758), .W4TO27(6161), .W4TO28(15846), .W4TO29(1104), .W4TO30(5098), .W4TO31(-12249), .W4TO32(-6429), .W4TO33(-830), .W4TO34(-1515), .W4TO35(4252), .W4TO36(-19503), .W4TO37(-1030), .W4TO38(20060), .W4TO39(5396), .W4TO40(-24116), .W4TO41(9069), .W4TO42(-4408), .W4TO43(-846), .W4TO44(18302), .W4TO45(-17468), .W4TO46(-11309), .W4TO47(-6685), .W4TO48(-11048), .W4TO49(12689), .W4TO50(253), .W4TO51(1262), .W4TO52(-72), .W4TO53(18178), .W4TO54(-181), .W4TO55(-9221), .W4TO56(-5824), .W4TO57(-1575), .W4TO58(-14518), .W4TO59(-1271), .W4TO60(-9482), .W4TO61(2807), .W4TO62(3067), .W4TO63(-12377), .W4TO64(-3052), .W4TO65(14330), .W4TO66(572), .W4TO67(-7779), .W4TO68(15590), .W4TO69(9580), .W4TO70(-746), .W4TO71(9375), .W4TO72(-4153), .W4TO73(-3082), .W4TO74(5842), .W4TO75(-19019), .W4TO76(10776), .W4TO77(-6075), .W4TO78(-3935), .W4TO79(-9280), .W4TO80(347), .W4TO81(18877), .W4TO82(-10549), .W4TO83(15974), .W4TO84(-24565), .W4TO85(18678), .W4TO86(-4297), .W4TO87(16649), .W4TO88(-13153), .W4TO89(-18857), .W4TO90(4261), .W4TO91(-3262), .W4TO92(17427), .W4TO93(14804), .W4TO94(8477), .W4TO95(-11182), .W4TO96(14854), .W4TO97(-8425), .W4TO98(-22322), .W4TO99(-1291), .W5TO0(-7265), .W5TO1(-1971), .W5TO2(1332), .W5TO3(-3078), .W5TO4(-23641), .W5TO5(-348), .W5TO6(8496), .W5TO7(12122), .W5TO8(-4868), .W5TO9(13747), .W5TO10(15840), .W5TO11(10611), .W5TO12(8654), .W5TO13(179), .W5TO14(4119), .W5TO15(-1980), .W5TO16(17305), .W5TO17(-6012), .W5TO18(6201), .W5TO19(1901), .W5TO20(3360), .W5TO21(313), .W5TO22(-4634), .W5TO23(-8066), .W5TO24(-60), .W5TO25(-10234), .W5TO26(-12446), .W5TO27(-500), .W5TO28(-17795), .W5TO29(-29035), .W5TO30(-19115), .W5TO31(-7933), .W5TO32(-11308), .W5TO33(3287), .W5TO34(-11020), .W5TO35(8515), .W5TO36(-17399), .W5TO37(3678), .W5TO38(-2113), .W5TO39(-10194), .W5TO40(10345), .W5TO41(-17917), .W5TO42(2684), .W5TO43(-5130), .W5TO44(-11586), .W5TO45(-5832), .W5TO46(-555), .W5TO47(12001), .W5TO48(6321), .W5TO49(-4290), .W5TO50(-15565), .W5TO51(13926), .W5TO52(10195), .W5TO53(13875), .W5TO54(-3547), .W5TO55(13832), .W5TO56(-5695), .W5TO57(941), .W5TO58(5807), .W5TO59(-5571), .W5TO60(1425), .W5TO61(22807), .W5TO62(9747), .W5TO63(-3430), .W5TO64(841), .W5TO65(13862), .W5TO66(-14809), .W5TO67(14309), .W5TO68(11974), .W5TO69(8190), .W5TO70(-15655), .W5TO71(-3038), .W5TO72(9909), .W5TO73(-14427), .W5TO74(241), .W5TO75(-7176), .W5TO76(6014), .W5TO77(13109), .W5TO78(-3626), .W5TO79(23612), .W5TO80(6632), .W5TO81(-5693), .W5TO82(11890), .W5TO83(2117), .W5TO84(-14100), .W5TO85(-10021), .W5TO86(-6946), .W5TO87(-14891), .W5TO88(-6539), .W5TO89(19612), .W5TO90(18208), .W5TO91(-7482), .W5TO92(-14270), .W5TO93(-14310), .W5TO94(-13006), .W5TO95(5314), .W5TO96(16918), .W5TO97(-13124), .W5TO98(-3635), .W5TO99(15727), .W6TO0(1963), .W6TO1(-5650), .W6TO2(-17626), .W6TO3(-9894), .W6TO4(-1412), .W6TO5(5537), .W6TO6(11379), .W6TO7(11338), .W6TO8(-5757), .W6TO9(-16250), .W6TO10(-12309), .W6TO11(-6657), .W6TO12(9591), .W6TO13(-7534), .W6TO14(-3673), .W6TO15(2944), .W6TO16(-1932), .W6TO17(1996), .W6TO18(-6632), .W6TO19(-16295), .W6TO20(-14535), .W6TO21(6771), .W6TO22(-2347), .W6TO23(-12286), .W6TO24(14248), .W6TO25(5280), .W6TO26(-7872), .W6TO27(-3358), .W6TO28(-6860), .W6TO29(13201), .W6TO30(-16704), .W6TO31(-18409), .W6TO32(64), .W6TO33(-435), .W6TO34(3543), .W6TO35(-3034), .W6TO36(16213), .W6TO37(-172), .W6TO38(6100), .W6TO39(-6279), .W6TO40(2066), .W6TO41(8192), .W6TO42(-18392), .W6TO43(-6727), .W6TO44(6014), .W6TO45(6088), .W6TO46(785), .W6TO47(8966), .W6TO48(-8084), .W6TO49(-10780), .W6TO50(-10665), .W6TO51(14551), .W6TO52(5594), .W6TO53(-3260), .W6TO54(-15527), .W6TO55(-18954), .W6TO56(-16546), .W6TO57(-11389), .W6TO58(-18310), .W6TO59(2948), .W6TO60(-13579), .W6TO61(-17400), .W6TO62(-8673), .W6TO63(-4025), .W6TO64(18383), .W6TO65(7663), .W6TO66(6011), .W6TO67(-11111), .W6TO68(13707), .W6TO69(-7294), .W6TO70(-9326), .W6TO71(-5244), .W6TO72(11984), .W6TO73(10545), .W6TO74(-18812), .W6TO75(14118), .W6TO76(-11161), .W6TO77(13795), .W6TO78(18009), .W6TO79(-4462), .W6TO80(-20718), .W6TO81(134), .W6TO82(-1962), .W6TO83(18238), .W6TO84(857), .W6TO85(10738), .W6TO86(11157), .W6TO87(14318), .W6TO88(10605), .W6TO89(-11885), .W6TO90(-12561), .W6TO91(1299), .W6TO92(9385), .W6TO93(6804), .W6TO94(-7282), .W6TO95(4461), .W6TO96(18389), .W6TO97(8733), .W6TO98(-19179), .W6TO99(17187), .W7TO0(5973), .W7TO1(-15166), .W7TO2(-17180), .W7TO3(8223), .W7TO4(11135), .W7TO5(-7241), .W7TO6(-4705), .W7TO7(9931), .W7TO8(-992), .W7TO9(-7618), .W7TO10(-5805), .W7TO11(-6569), .W7TO12(10636), .W7TO13(14181), .W7TO14(-3137), .W7TO15(-13364), .W7TO16(7971), .W7TO17(-15244), .W7TO18(8049), .W7TO19(13125), .W7TO20(-12643), .W7TO21(-11948), .W7TO22(-15655), .W7TO23(-17975), .W7TO24(-8481), .W7TO25(9160), .W7TO26(-4173), .W7TO27(-14613), .W7TO28(10898), .W7TO29(5478), .W7TO30(-15167), .W7TO31(17763), .W7TO32(13709), .W7TO33(-2638), .W7TO34(-9972), .W7TO35(-6587), .W7TO36(8843), .W7TO37(13914), .W7TO38(-2351), .W7TO39(-1899), .W7TO40(1946), .W7TO41(2371), .W7TO42(1664), .W7TO43(-1248), .W7TO44(12613), .W7TO45(3019), .W7TO46(5594), .W7TO47(10505), .W7TO48(3647), .W7TO49(-6487), .W7TO50(3454), .W7TO51(2011), .W7TO52(12119), .W7TO53(-13485), .W7TO54(-18740), .W7TO55(-15595), .W7TO56(-3577), .W7TO57(-8200), .W7TO58(4621), .W7TO59(6512), .W7TO60(3607), .W7TO61(15771), .W7TO62(-13323), .W7TO63(15678), .W7TO64(-7592), .W7TO65(-4778), .W7TO66(-2225), .W7TO67(-98), .W7TO68(7257), .W7TO69(1929), .W7TO70(-13855), .W7TO71(18791), .W7TO72(-1335), .W7TO73(2969), .W7TO74(13081), .W7TO75(1605), .W7TO76(-19231), .W7TO77(-12946), .W7TO78(-133), .W7TO79(-13067), .W7TO80(5344), .W7TO81(-15973), .W7TO82(-13437), .W7TO83(854), .W7TO84(14633), .W7TO85(-18131), .W7TO86(-6151), .W7TO87(-6253), .W7TO88(-10141), .W7TO89(19214), .W7TO90(3293), .W7TO91(7885), .W7TO92(17820), .W7TO93(4909), .W7TO94(17193), .W7TO95(-11732), .W7TO96(11239), .W7TO97(-4610), .W7TO98(-10632), .W7TO99(-13595), .W8TO0(8881), .W8TO1(-15936), .W8TO2(2625), .W8TO3(12452), .W8TO4(-14810), .W8TO5(-15104), .W8TO6(-9109), .W8TO7(-9886), .W8TO8(-2623), .W8TO9(9434), .W8TO10(-18890), .W8TO11(-10048), .W8TO12(-16896), .W8TO13(-8274), .W8TO14(15921), .W8TO15(11420), .W8TO16(-6901), .W8TO17(345), .W8TO18(-17611), .W8TO19(12739), .W8TO20(-6448), .W8TO21(-17334), .W8TO22(6320), .W8TO23(12391), .W8TO24(-9510), .W8TO25(10209), .W8TO26(8099), .W8TO27(-680), .W8TO28(-9397), .W8TO29(5496), .W8TO30(16662), .W8TO31(5599), .W8TO32(-13217), .W8TO33(-10735), .W8TO34(6767), .W8TO35(4540), .W8TO36(7323), .W8TO37(2582), .W8TO38(7625), .W8TO39(-14015), .W8TO40(11813), .W8TO41(-2758), .W8TO42(-17075), .W8TO43(-3177), .W8TO44(15127), .W8TO45(-11868), .W8TO46(4945), .W8TO47(17404), .W8TO48(9193), .W8TO49(-15501), .W8TO50(-5866), .W8TO51(-11709), .W8TO52(-5405), .W8TO53(18482), .W8TO54(-17729), .W8TO55(-3669), .W8TO56(2736), .W8TO57(-11809), .W8TO58(17591), .W8TO59(12759), .W8TO60(8084), .W8TO61(17477), .W8TO62(-11695), .W8TO63(-16738), .W8TO64(-8637), .W8TO65(12764), .W8TO66(2082), .W8TO67(-5525), .W8TO68(-16917), .W8TO69(-1025), .W8TO70(10970), .W8TO71(11142), .W8TO72(-9744), .W8TO73(-1577), .W8TO74(-7300), .W8TO75(-2515), .W8TO76(11673), .W8TO77(-4480), .W8TO78(1682), .W8TO79(-3211), .W8TO80(-11820), .W8TO81(10995), .W8TO82(-12517), .W8TO83(-5752), .W8TO84(11191), .W8TO85(13144), .W8TO86(-16798), .W8TO87(-481), .W8TO88(-10524), .W8TO89(-9659), .W8TO90(12531), .W8TO91(6576), .W8TO92(-10688), .W8TO93(-5864), .W8TO94(18422), .W8TO95(3499), .W8TO96(17579), .W8TO97(-18822), .W8TO98(1133), .W8TO99(18567), .W9TO0(-14600), .W9TO1(9244), .W9TO2(4426), .W9TO3(-10811), .W9TO4(-3103), .W9TO5(-14160), .W9TO6(12563), .W9TO7(6483), .W9TO8(13689), .W9TO9(2739), .W9TO10(976), .W9TO11(3380), .W9TO12(-5824), .W9TO13(-3962), .W9TO14(-13311), .W9TO15(9351), .W9TO16(-7189), .W9TO17(-5099), .W9TO18(-2656), .W9TO19(-10727), .W9TO20(-12416), .W9TO21(860), .W9TO22(-11317), .W9TO23(-11906), .W9TO24(7456), .W9TO25(-13130), .W9TO26(8153), .W9TO27(-117), .W9TO28(16685), .W9TO29(-13804), .W9TO30(-11912), .W9TO31(2391), .W9TO32(-256), .W9TO33(-7230), .W9TO34(9097), .W9TO35(-3337), .W9TO36(5332), .W9TO37(-6436), .W9TO38(2201), .W9TO39(-19120), .W9TO40(-11633), .W9TO41(-5067), .W9TO42(-3776), .W9TO43(8415), .W9TO44(-19030), .W9TO45(-11015), .W9TO46(14880), .W9TO47(-7100), .W9TO48(-10547), .W9TO49(-16935), .W9TO50(3639), .W9TO51(16039), .W9TO52(17234), .W9TO53(11543), .W9TO54(-7413), .W9TO55(-718), .W9TO56(-12491), .W9TO57(18948), .W9TO58(4818), .W9TO59(3284), .W9TO60(-13304), .W9TO61(-9487), .W9TO62(-13356), .W9TO63(-4887), .W9TO64(11250), .W9TO65(-3103), .W9TO66(-2210), .W9TO67(10486), .W9TO68(15418), .W9TO69(-2450), .W9TO70(-7319), .W9TO71(8052), .W9TO72(11536), .W9TO73(-1419), .W9TO74(-13128), .W9TO75(-9247), .W9TO76(-7898), .W9TO77(-11322), .W9TO78(-10929), .W9TO79(12141), .W9TO80(11442), .W9TO81(3131), .W9TO82(18075), .W9TO83(18144), .W9TO84(-15136), .W9TO85(-17159), .W9TO86(541), .W9TO87(-16510), .W9TO88(1006), .W9TO89(16345), .W9TO90(4270), .W9TO91(13901), .W9TO92(-5644), .W9TO93(-14063), .W9TO94(-18139), .W9TO95(-7647), .W9TO96(7367), .W9TO97(-15954), .W9TO98(-3899), .W9TO99(9305), .W10TO0(-18368), .W10TO1(7852), .W10TO2(2262), .W10TO3(-16804), .W10TO4(445), .W10TO5(7368), .W10TO6(-16809), .W10TO7(1895), .W10TO8(-1090), .W10TO9(17165), .W10TO10(-19925), .W10TO11(-1044), .W10TO12(18307), .W10TO13(-4200), .W10TO14(12370), .W10TO15(7419), .W10TO16(-12310), .W10TO17(3180), .W10TO18(15344), .W10TO19(-6507), .W10TO20(3384), .W10TO21(-13771), .W10TO22(-466), .W10TO23(3477), .W10TO24(25807), .W10TO25(-15589), .W10TO26(-14909), .W10TO27(-2770), .W10TO28(2948), .W10TO29(6944), .W10TO30(9420), .W10TO31(59), .W10TO32(-12042), .W10TO33(10782), .W10TO34(-280), .W10TO35(-5348), .W10TO36(7733), .W10TO37(1416), .W10TO38(-2490), .W10TO39(-6004), .W10TO40(-701), .W10TO41(-16824), .W10TO42(-5160), .W10TO43(-3063), .W10TO44(2381), .W10TO45(13399), .W10TO46(-18723), .W10TO47(2839), .W10TO48(6564), .W10TO49(-10782), .W10TO50(-4244), .W10TO51(2909), .W10TO52(6372), .W10TO53(-3009), .W10TO54(2024), .W10TO55(5833), .W10TO56(2632), .W10TO57(5266), .W10TO58(7834), .W10TO59(-4627), .W10TO60(-25167), .W10TO61(-6587), .W10TO62(-10911), .W10TO63(15146), .W10TO64(17691), .W10TO65(-15919), .W10TO66(-1538), .W10TO67(7142), .W10TO68(-5189), .W10TO69(5335), .W10TO70(13215), .W10TO71(-13742), .W10TO72(9413), .W10TO73(-10631), .W10TO74(-8877), .W10TO75(-18974), .W10TO76(2044), .W10TO77(-15936), .W10TO78(-5029), .W10TO79(-9168), .W10TO80(7551), .W10TO81(-12509), .W10TO82(14221), .W10TO83(9214), .W10TO84(-11631), .W10TO85(12726), .W10TO86(9441), .W10TO87(679), .W10TO88(-12688), .W10TO89(-8963), .W10TO90(-10998), .W10TO91(4601), .W10TO92(-2932), .W10TO93(-6498), .W10TO94(7482), .W10TO95(5911), .W10TO96(18175), .W10TO97(12335), .W10TO98(-16628), .W10TO99(-3767), .W11TO0(-288), .W11TO1(-9604), .W11TO2(11193), .W11TO3(4788), .W11TO4(14736), .W11TO5(8052), .W11TO6(2810), .W11TO7(10095), .W11TO8(-11229), .W11TO9(2177), .W11TO10(14350), .W11TO11(13574), .W11TO12(14170), .W11TO13(-1103), .W11TO14(13184), .W11TO15(-4777), .W11TO16(8964), .W11TO17(-6277), .W11TO18(-10904), .W11TO19(-8308), .W11TO20(-14455), .W11TO21(5879), .W11TO22(-13734), .W11TO23(8295), .W11TO24(-4696), .W11TO25(-11569), .W11TO26(-18419), .W11TO27(-15724), .W11TO28(3524), .W11TO29(-1951), .W11TO30(18111), .W11TO31(8300), .W11TO32(4494), .W11TO33(12658), .W11TO34(-15124), .W11TO35(5990), .W11TO36(-7808), .W11TO37(-497), .W11TO38(18709), .W11TO39(6805), .W11TO40(-2654), .W11TO41(6939), .W11TO42(6091), .W11TO43(6134), .W11TO44(15317), .W11TO45(-22439), .W11TO46(-11326), .W11TO47(5109), .W11TO48(-14055), .W11TO49(5090), .W11TO50(13809), .W11TO51(-2451), .W11TO52(9616), .W11TO53(-6199), .W11TO54(514), .W11TO55(16072), .W11TO56(-4329), .W11TO57(-6523), .W11TO58(5782), .W11TO59(8556), .W11TO60(15825), .W11TO61(-10426), .W11TO62(-14732), .W11TO63(-10929), .W11TO64(17534), .W11TO65(-8590), .W11TO66(-18276), .W11TO67(10424), .W11TO68(1105), .W11TO69(21124), .W11TO70(1933), .W11TO71(12372), .W11TO72(8136), .W11TO73(-10393), .W11TO74(-8323), .W11TO75(2179), .W11TO76(-1225), .W11TO77(8720), .W11TO78(998), .W11TO79(169), .W11TO80(-4989), .W11TO81(15158), .W11TO82(-10911), .W11TO83(1079), .W11TO84(5343), .W11TO85(1642), .W11TO86(-15033), .W11TO87(12477), .W11TO88(-16427), .W11TO89(-8162), .W11TO90(-1368), .W11TO91(-10907), .W11TO92(-107), .W11TO93(324), .W11TO94(-21440), .W11TO95(-477), .W11TO96(-4558), .W11TO97(-5241), .W11TO98(6993), .W11TO99(11860), .W12TO0(-11237), .W12TO1(-6705), .W12TO2(6104), .W12TO3(4275), .W12TO4(3801), .W12TO5(-16094), .W12TO6(-17694), .W12TO7(21541), .W12TO8(17512), .W12TO9(11621), .W12TO10(13758), .W12TO11(-9225), .W12TO12(15091), .W12TO13(4513), .W12TO14(-1324), .W12TO15(-2487), .W12TO16(706), .W12TO17(-3873), .W12TO18(-3708), .W12TO19(8263), .W12TO20(14347), .W12TO21(19247), .W12TO22(-3328), .W12TO23(5853), .W12TO24(-6327), .W12TO25(-7284), .W12TO26(6815), .W12TO27(-6219), .W12TO28(-15535), .W12TO29(1817), .W12TO30(-21466), .W12TO31(-19798), .W12TO32(3592), .W12TO33(-15832), .W12TO34(7202), .W12TO35(-16219), .W12TO36(-8047), .W12TO37(13205), .W12TO38(477), .W12TO39(4925), .W12TO40(-13917), .W12TO41(-12846), .W12TO42(-7568), .W12TO43(-18400), .W12TO44(11367), .W12TO45(-9963), .W12TO46(5050), .W12TO47(13577), .W12TO48(-21429), .W12TO49(-4030), .W12TO50(4702), .W12TO51(550), .W12TO52(15101), .W12TO53(2409), .W12TO54(-6524), .W12TO55(6353), .W12TO56(13411), .W12TO57(5800), .W12TO58(2913), .W12TO59(16999), .W12TO60(945), .W12TO61(16432), .W12TO62(-7822), .W12TO63(-13125), .W12TO64(-6788), .W12TO65(9111), .W12TO66(195), .W12TO67(510), .W12TO68(19959), .W12TO69(19189), .W12TO70(-18118), .W12TO71(-10968), .W12TO72(-9061), .W12TO73(-21553), .W12TO74(-12688), .W12TO75(17496), .W12TO76(3148), .W12TO77(-16968), .W12TO78(2714), .W12TO79(18587), .W12TO80(1269), .W12TO81(16072), .W12TO82(-20279), .W12TO83(-1820), .W12TO84(-17021), .W12TO85(-6315), .W12TO86(2297), .W12TO87(-4585), .W12TO88(-4816), .W12TO89(16745), .W12TO90(2948), .W12TO91(2496), .W12TO92(19025), .W12TO93(-13958), .W12TO94(-19815), .W12TO95(-21352), .W12TO96(17793), .W12TO97(3169), .W12TO98(2209), .W12TO99(-7843), .W13TO0(10323), .W13TO1(10609), .W13TO2(14468), .W13TO3(13661), .W13TO4(-5279), .W13TO5(9005), .W13TO6(-12383), .W13TO7(-10653), .W13TO8(4769), .W13TO9(12382), .W13TO10(5215), .W13TO11(14843), .W13TO12(7457), .W13TO13(12061), .W13TO14(1044), .W13TO15(7282), .W13TO16(13426), .W13TO17(19401), .W13TO18(-20267), .W13TO19(7371), .W13TO20(-1661), .W13TO21(1810), .W13TO22(4690), .W13TO23(-10258), .W13TO24(20869), .W13TO25(-13857), .W13TO26(9439), .W13TO27(12321), .W13TO28(-13515), .W13TO29(4227), .W13TO30(-11292), .W13TO31(9105), .W13TO32(-3064), .W13TO33(14190), .W13TO34(-3783), .W13TO35(5369), .W13TO36(11014), .W13TO37(19389), .W13TO38(2411), .W13TO39(-765), .W13TO40(-5469), .W13TO41(84), .W13TO42(-16166), .W13TO43(18366), .W13TO44(1831), .W13TO45(-5323), .W13TO46(18523), .W13TO47(-2788), .W13TO48(-13733), .W13TO49(6217), .W13TO50(11834), .W13TO51(-9051), .W13TO52(-10502), .W13TO53(-1797), .W13TO54(6574), .W13TO55(-2781), .W13TO56(1952), .W13TO57(-18069), .W13TO58(-13288), .W13TO59(6453), .W13TO60(-5397), .W13TO61(26448), .W13TO62(-13613), .W13TO63(-1702), .W13TO64(-13153), .W13TO65(-18751), .W13TO66(9643), .W13TO67(-11327), .W13TO68(10399), .W13TO69(-6072), .W13TO70(-8213), .W13TO71(-3403), .W13TO72(21260), .W13TO73(-3517), .W13TO74(-17626), .W13TO75(-5351), .W13TO76(-5281), .W13TO77(5925), .W13TO78(-894), .W13TO79(23306), .W13TO80(4932), .W13TO81(-8805), .W13TO82(-4213), .W13TO83(5314), .W13TO84(9421), .W13TO85(18972), .W13TO86(-16847), .W13TO87(7520), .W13TO88(6887), .W13TO89(15365), .W13TO90(-221), .W13TO91(3430), .W13TO92(10926), .W13TO93(-8221), .W13TO94(-14695), .W13TO95(-9713), .W13TO96(8953), .W13TO97(-17582), .W13TO98(-10751), .W13TO99(8804), .W14TO0(-17676), .W14TO1(4771), .W14TO2(2926), .W14TO3(-13873), .W14TO4(5113), .W14TO5(3071), .W14TO6(13830), .W14TO7(11920), .W14TO8(4140), .W14TO9(18714), .W14TO10(-22), .W14TO11(-6408), .W14TO12(6156), .W14TO13(11627), .W14TO14(7175), .W14TO15(-6201), .W14TO16(11065), .W14TO17(17833), .W14TO18(-14230), .W14TO19(11380), .W14TO20(-14680), .W14TO21(9448), .W14TO22(-11808), .W14TO23(15060), .W14TO24(15496), .W14TO25(-7569), .W14TO26(10808), .W14TO27(-17871), .W14TO28(-10181), .W14TO29(-7867), .W14TO30(-7173), .W14TO31(-974), .W14TO32(-3283), .W14TO33(3474), .W14TO34(-7490), .W14TO35(2522), .W14TO36(-17159), .W14TO37(4316), .W14TO38(-1434), .W14TO39(-8604), .W14TO40(-18379), .W14TO41(-11020), .W14TO42(-2607), .W14TO43(1117), .W14TO44(-811), .W14TO45(-7831), .W14TO46(10918), .W14TO47(794), .W14TO48(-746), .W14TO49(4665), .W14TO50(-10765), .W14TO51(5715), .W14TO52(15168), .W14TO53(-12089), .W14TO54(-4083), .W14TO55(11899), .W14TO56(19006), .W14TO57(12379), .W14TO58(11480), .W14TO59(7301), .W14TO60(-827), .W14TO61(2005), .W14TO62(-1551), .W14TO63(13823), .W14TO64(4146), .W14TO65(1786), .W14TO66(-17570), .W14TO67(6383), .W14TO68(-13207), .W14TO69(18773), .W14TO70(-12719), .W14TO71(1836), .W14TO72(-15568), .W14TO73(-11498), .W14TO74(-14876), .W14TO75(-13033), .W14TO76(-2561), .W14TO77(-3362), .W14TO78(-10178), .W14TO79(5343), .W14TO80(-313), .W14TO81(-11285), .W14TO82(7810), .W14TO83(-12892), .W14TO84(10299), .W14TO85(-5812), .W14TO86(-12350), .W14TO87(6463), .W14TO88(15562), .W14TO89(-54), .W14TO90(19482), .W14TO91(-16423), .W14TO92(-12851), .W14TO93(3919), .W14TO94(4144), .W14TO95(-18894), .W14TO96(10785), .W14TO97(8730), .W14TO98(10449), .W14TO99(18888), .W15TO0(-15239), .W15TO1(-663), .W15TO2(-3271), .W15TO3(9125), .W15TO4(13335), .W15TO5(-3545), .W15TO6(3037), .W15TO7(13340), .W15TO8(-18223), .W15TO9(15901), .W15TO10(-1297), .W15TO11(-6545), .W15TO12(9374), .W15TO13(15306), .W15TO14(-9575), .W15TO15(-8433), .W15TO16(15061), .W15TO17(1624), .W15TO18(-7213), .W15TO19(-10967), .W15TO20(-9721), .W15TO21(14720), .W15TO22(18448), .W15TO23(945), .W15TO24(10475), .W15TO25(3762), .W15TO26(-5518), .W15TO27(2881), .W15TO28(-14447), .W15TO29(5932), .W15TO30(3064), .W15TO31(-15248), .W15TO32(17872), .W15TO33(17451), .W15TO34(16368), .W15TO35(9570), .W15TO36(3577), .W15TO37(9064), .W15TO38(17320), .W15TO39(-17401), .W15TO40(2037), .W15TO41(-1326), .W15TO42(10709), .W15TO43(-1570), .W15TO44(14305), .W15TO45(1758), .W15TO46(-2063), .W15TO47(-15507), .W15TO48(-4775), .W15TO49(-10937), .W15TO50(8923), .W15TO51(-14786), .W15TO52(13003), .W15TO53(-4971), .W15TO54(11448), .W15TO55(19066), .W15TO56(-14054), .W15TO57(-2197), .W15TO58(16761), .W15TO59(-5780), .W15TO60(-16791), .W15TO61(11933), .W15TO62(6356), .W15TO63(-8526), .W15TO64(-17549), .W15TO65(-9541), .W15TO66(16027), .W15TO67(12951), .W15TO68(14110), .W15TO69(-540), .W15TO70(14299), .W15TO71(14746), .W15TO72(9257), .W15TO73(-3776), .W15TO74(2618), .W15TO75(-16990), .W15TO76(-1261), .W15TO77(-9257), .W15TO78(-18302), .W15TO79(-8216), .W15TO80(-11677), .W15TO81(17318), .W15TO82(13784), .W15TO83(15995), .W15TO84(9959), .W15TO85(-12406), .W15TO86(-3078), .W15TO87(8046), .W15TO88(-4829), .W15TO89(-6687), .W15TO90(-15085), .W15TO91(-517), .W15TO92(-10526), .W15TO93(-15067), .W15TO94(-9671), .W15TO95(6593), .W15TO96(-10603), .W15TO97(-13280), .W15TO98(-1242), .W15TO99(-2720), .W16TO0(-1569), .W16TO1(-5475), .W16TO2(-18955), .W16TO3(2518), .W16TO4(-3552), .W16TO5(7408), .W16TO6(16760), .W16TO7(-5050), .W16TO8(12253), .W16TO9(-12246), .W16TO10(9315), .W16TO11(-16183), .W16TO12(4309), .W16TO13(-12483), .W16TO14(-14731), .W16TO15(-3823), .W16TO16(-11047), .W16TO17(-12777), .W16TO18(13638), .W16TO19(12126), .W16TO20(16401), .W16TO21(-13847), .W16TO22(18229), .W16TO23(17147), .W16TO24(13966), .W16TO25(-10730), .W16TO26(4684), .W16TO27(7888), .W16TO28(-800), .W16TO29(15142), .W16TO30(12517), .W16TO31(7042), .W16TO32(-7204), .W16TO33(-13593), .W16TO34(40), .W16TO35(4532), .W16TO36(13393), .W16TO37(-3478), .W16TO38(-17637), .W16TO39(5930), .W16TO40(-9245), .W16TO41(7758), .W16TO42(-4800), .W16TO43(923), .W16TO44(17363), .W16TO45(-6040), .W16TO46(17958), .W16TO47(-2512), .W16TO48(12466), .W16TO49(18055), .W16TO50(18627), .W16TO51(-16419), .W16TO52(16825), .W16TO53(2615), .W16TO54(10479), .W16TO55(4251), .W16TO56(11181), .W16TO57(-13649), .W16TO58(14525), .W16TO59(-15178), .W16TO60(-4056), .W16TO61(1598), .W16TO62(-8363), .W16TO63(-13982), .W16TO64(5533), .W16TO65(8250), .W16TO66(11962), .W16TO67(15277), .W16TO68(13243), .W16TO69(5737), .W16TO70(2830), .W16TO71(7828), .W16TO72(-14992), .W16TO73(-994), .W16TO74(-12074), .W16TO75(4331), .W16TO76(-13169), .W16TO77(-16741), .W16TO78(16596), .W16TO79(7483), .W16TO80(-2855), .W16TO81(-2436), .W16TO82(-4451), .W16TO83(-1613), .W16TO84(12649), .W16TO85(-1317), .W16TO86(14678), .W16TO87(15811), .W16TO88(-17449), .W16TO89(2034), .W16TO90(452), .W16TO91(-14745), .W16TO92(-9791), .W16TO93(11021), .W16TO94(4101), .W16TO95(13421), .W16TO96(-1382), .W16TO97(11660), .W16TO98(-11207), .W16TO99(18426), .W17TO0(2173), .W17TO1(15911), .W17TO2(-15223), .W17TO3(14316), .W17TO4(-1907), .W17TO5(-13942), .W17TO6(5288), .W17TO7(-20752), .W17TO8(10332), .W17TO9(13405), .W17TO10(-9186), .W17TO11(-17787), .W17TO12(-5062), .W17TO13(7932), .W17TO14(-10229), .W17TO15(-17328), .W17TO16(-3634), .W17TO17(17993), .W17TO18(-3184), .W17TO19(-7251), .W17TO20(16310), .W17TO21(-860), .W17TO22(20009), .W17TO23(13862), .W17TO24(12582), .W17TO25(-638), .W17TO26(-4056), .W17TO27(-2188), .W17TO28(94), .W17TO29(7303), .W17TO30(-2357), .W17TO31(-21197), .W17TO32(9237), .W17TO33(10029), .W17TO34(-11549), .W17TO35(3805), .W17TO36(2402), .W17TO37(-11898), .W17TO38(-8644), .W17TO39(-12673), .W17TO40(16164), .W17TO41(3943), .W17TO42(16423), .W17TO43(-1010), .W17TO44(10082), .W17TO45(13323), .W17TO46(4229), .W17TO47(3115), .W17TO48(14758), .W17TO49(584), .W17TO50(-6026), .W17TO51(11139), .W17TO52(12931), .W17TO53(11246), .W17TO54(-15636), .W17TO55(3019), .W17TO56(-12073), .W17TO57(16035), .W17TO58(-284), .W17TO59(466), .W17TO60(-11650), .W17TO61(-11865), .W17TO62(11759), .W17TO63(-5109), .W17TO64(7342), .W17TO65(14924), .W17TO66(3342), .W17TO67(-11657), .W17TO68(17139), .W17TO69(17160), .W17TO70(4176), .W17TO71(-15841), .W17TO72(14966), .W17TO73(-12393), .W17TO74(15668), .W17TO75(-6954), .W17TO76(-8940), .W17TO77(11025), .W17TO78(1315), .W17TO79(4452), .W17TO80(-5577), .W17TO81(-13002), .W17TO82(-11035), .W17TO83(-1813), .W17TO84(-7778), .W17TO85(-13084), .W17TO86(-8078), .W17TO87(4230), .W17TO88(-5179), .W17TO89(-84), .W17TO90(-11417), .W17TO91(3727), .W17TO92(6799), .W17TO93(3058), .W17TO94(8), .W17TO95(7503), .W17TO96(-9162), .W17TO97(4473), .W17TO98(-14253), .W17TO99(-12304), .W18TO0(-4110), .W18TO1(2421), .W18TO2(10615), .W18TO3(-10856), .W18TO4(15997), .W18TO5(4320), .W18TO6(12868), .W18TO7(-3179), .W18TO8(1346), .W18TO9(-5950), .W18TO10(3700), .W18TO11(15779), .W18TO12(10741), .W18TO13(-6244), .W18TO14(-18211), .W18TO15(-11631), .W18TO16(12891), .W18TO17(16368), .W18TO18(9310), .W18TO19(-13373), .W18TO20(9992), .W18TO21(14905), .W18TO22(-8492), .W18TO23(-11226), .W18TO24(377), .W18TO25(-12106), .W18TO26(-987), .W18TO27(-8219), .W18TO28(-17322), .W18TO29(-10961), .W18TO30(20030), .W18TO31(-17249), .W18TO32(-4049), .W18TO33(1975), .W18TO34(-11200), .W18TO35(17281), .W18TO36(8203), .W18TO37(13217), .W18TO38(5132), .W18TO39(3960), .W18TO40(-12142), .W18TO41(6944), .W18TO42(-15830), .W18TO43(6304), .W18TO44(-12121), .W18TO45(7464), .W18TO46(2452), .W18TO47(-1131), .W18TO48(1765), .W18TO49(7295), .W18TO50(2993), .W18TO51(-6242), .W18TO52(10633), .W18TO53(-16927), .W18TO54(16765), .W18TO55(6768), .W18TO56(11758), .W18TO57(-1710), .W18TO58(-11300), .W18TO59(6101), .W18TO60(3389), .W18TO61(-3131), .W18TO62(3756), .W18TO63(11049), .W18TO64(-8903), .W18TO65(17453), .W18TO66(-6233), .W18TO67(-21696), .W18TO68(-8140), .W18TO69(-35), .W18TO70(14691), .W18TO71(-12313), .W18TO72(-7735), .W18TO73(-20109), .W18TO74(-18243), .W18TO75(-4047), .W18TO76(-4636), .W18TO77(-9277), .W18TO78(-17925), .W18TO79(-9970), .W18TO80(4883), .W18TO81(-5938), .W18TO82(14329), .W18TO83(7654), .W18TO84(19707), .W18TO85(-9896), .W18TO86(6709), .W18TO87(13546), .W18TO88(-1591), .W18TO89(9869), .W18TO90(1592), .W18TO91(-5538), .W18TO92(19153), .W18TO93(-19211), .W18TO94(608), .W18TO95(-22834), .W18TO96(-3220), .W18TO97(6125), .W18TO98(12491), .W18TO99(4785), .W19TO0(-14329), .W19TO1(-16253), .W19TO2(-8778), .W19TO3(16013), .W19TO4(-8564), .W19TO5(7108), .W19TO6(-8680), .W19TO7(-13138), .W19TO8(5244), .W19TO9(-4899), .W19TO10(-15158), .W19TO11(7395), .W19TO12(-1135), .W19TO13(-9961), .W19TO14(-4166), .W19TO15(7085), .W19TO16(3093), .W19TO17(-4195), .W19TO18(-1371), .W19TO19(-7083), .W19TO20(7976), .W19TO21(350), .W19TO22(-3431), .W19TO23(-4478), .W19TO24(-6758), .W19TO25(-4088), .W19TO26(-23075), .W19TO27(-10851), .W19TO28(-10908), .W19TO29(-5374), .W19TO30(-14451), .W19TO31(-1471), .W19TO32(11814), .W19TO33(-7280), .W19TO34(-19083), .W19TO35(2463), .W19TO36(12175), .W19TO37(-6332), .W19TO38(7005), .W19TO39(10739), .W19TO40(-8443), .W19TO41(-10054), .W19TO42(12751), .W19TO43(-12307), .W19TO44(10534), .W19TO45(-15614), .W19TO46(13708), .W19TO47(1582), .W19TO48(10795), .W19TO49(11221), .W19TO50(5162), .W19TO51(-11816), .W19TO52(-8201), .W19TO53(6153), .W19TO54(11222), .W19TO55(15903), .W19TO56(-3145), .W19TO57(3376), .W19TO58(-21341), .W19TO59(-2275), .W19TO60(22093), .W19TO61(-5707), .W19TO62(-15975), .W19TO63(-8017), .W19TO64(3263), .W19TO65(19322), .W19TO66(-3094), .W19TO67(-14065), .W19TO68(11434), .W19TO69(4965), .W19TO70(-15445), .W19TO71(-5018), .W19TO72(7648), .W19TO73(-14948), .W19TO74(-18495), .W19TO75(-11133), .W19TO76(5841), .W19TO77(-15326), .W19TO78(-1722), .W19TO79(9205), .W19TO80(5746), .W19TO81(2431), .W19TO82(5318), .W19TO83(-16852), .W19TO84(15977), .W19TO85(10806), .W19TO86(20213), .W19TO87(-9985), .W19TO88(13849), .W19TO89(9623), .W19TO90(13127), .W19TO91(-9540), .W19TO92(5790), .W19TO93(-4530), .W19TO94(7965), .W19TO95(-10631), .W19TO96(-7978), .W19TO97(14733), .W19TO98(17734), .W19TO99(6941), .W20TO0(2661), .W20TO1(5012), .W20TO2(-8063), .W20TO3(6827), .W20TO4(-12290), .W20TO5(-2795), .W20TO6(5520), .W20TO7(-16047), .W20TO8(-17701), .W20TO9(-12154), .W20TO10(16348), .W20TO11(-8795), .W20TO12(-4550), .W20TO13(14634), .W20TO14(18172), .W20TO15(17684), .W20TO16(-20716), .W20TO17(17055), .W20TO18(17124), .W20TO19(17969), .W20TO20(-24260), .W20TO21(-9313), .W20TO22(-2767), .W20TO23(-12187), .W20TO24(-11995), .W20TO25(2637), .W20TO26(-4171), .W20TO27(-14271), .W20TO28(-2806), .W20TO29(-8947), .W20TO30(97), .W20TO31(-5051), .W20TO32(3204), .W20TO33(2721), .W20TO34(13508), .W20TO35(-1196), .W20TO36(-14958), .W20TO37(10846), .W20TO38(7493), .W20TO39(-7581), .W20TO40(-2511), .W20TO41(1712), .W20TO42(-17075), .W20TO43(13995), .W20TO44(-15047), .W20TO45(-20763), .W20TO46(-14741), .W20TO47(27549), .W20TO48(-18876), .W20TO49(-12417), .W20TO50(-13613), .W20TO51(-10189), .W20TO52(-14268), .W20TO53(5072), .W20TO54(4669), .W20TO55(1380), .W20TO56(-8342), .W20TO57(6175), .W20TO58(4166), .W20TO59(-20517), .W20TO60(7395), .W20TO61(-3698), .W20TO62(-3294), .W20TO63(92), .W20TO64(-13765), .W20TO65(5329), .W20TO66(-7542), .W20TO67(-11687), .W20TO68(-11457), .W20TO69(1927), .W20TO70(2603), .W20TO71(-8435), .W20TO72(16105), .W20TO73(11426), .W20TO74(-13526), .W20TO75(-8940), .W20TO76(10610), .W20TO77(18914), .W20TO78(11495), .W20TO79(-6124), .W20TO80(-12427), .W20TO81(13354), .W20TO82(189), .W20TO83(-7565), .W20TO84(2705), .W20TO85(-3765), .W20TO86(8022), .W20TO87(-22868), .W20TO88(-4496), .W20TO89(6292), .W20TO90(13015), .W20TO91(14438), .W20TO92(305), .W20TO93(1664), .W20TO94(-2970), .W20TO95(8070), .W20TO96(5385), .W20TO97(-3284), .W20TO98(7041), .W20TO99(3971), .W21TO0(-11909), .W21TO1(4995), .W21TO2(6525), .W21TO3(-18752), .W21TO4(11174), .W21TO5(-33567), .W21TO6(-3856), .W21TO7(-7967), .W21TO8(-5853), .W21TO9(4888), .W21TO10(-9403), .W21TO11(20037), .W21TO12(4207), .W21TO13(14128), .W21TO14(-245), .W21TO15(21034), .W21TO16(-4478), .W21TO17(-10337), .W21TO18(-15717), .W21TO19(1530), .W21TO20(-22063), .W21TO21(12512), .W21TO22(17257), .W21TO23(9530), .W21TO24(17038), .W21TO25(14967), .W21TO26(-18310), .W21TO27(-5791), .W21TO28(-9319), .W21TO29(11988), .W21TO30(-1715), .W21TO31(-7802), .W21TO32(-2888), .W21TO33(-25191), .W21TO34(9966), .W21TO35(1840), .W21TO36(-18623), .W21TO37(18980), .W21TO38(9136), .W21TO39(-4680), .W21TO40(12150), .W21TO41(10222), .W21TO42(-9360), .W21TO43(-3223), .W21TO44(-17557), .W21TO45(7411), .W21TO46(-9974), .W21TO47(24547), .W21TO48(-15187), .W21TO49(-9366), .W21TO50(16254), .W21TO51(8554), .W21TO52(9575), .W21TO53(-25324), .W21TO54(-19165), .W21TO55(-3134), .W21TO56(-13181), .W21TO57(-2684), .W21TO58(13783), .W21TO59(-4045), .W21TO60(-584), .W21TO61(13035), .W21TO62(-15525), .W21TO63(17536), .W21TO64(-3268), .W21TO65(-7932), .W21TO66(10168), .W21TO67(-7736), .W21TO68(11391), .W21TO69(13821), .W21TO70(16312), .W21TO71(21166), .W21TO72(-6045), .W21TO73(13009), .W21TO74(11834), .W21TO75(7244), .W21TO76(-17337), .W21TO77(-10990), .W21TO78(-3503), .W21TO79(-17292), .W21TO80(14732), .W21TO81(217), .W21TO82(944), .W21TO83(-3063), .W21TO84(2877), .W21TO85(-4384), .W21TO86(8363), .W21TO87(5930), .W21TO88(-62), .W21TO89(6775), .W21TO90(2325), .W21TO91(-3020), .W21TO92(-349), .W21TO93(252), .W21TO94(1017), .W21TO95(1712), .W21TO96(-7303), .W21TO97(-12950), .W21TO98(11020), .W21TO99(13621), .W22TO0(-6587), .W22TO1(5746), .W22TO2(-12384), .W22TO3(-19284), .W22TO4(-15253), .W22TO5(-13622), .W22TO6(6524), .W22TO7(-10494), .W22TO8(-5329), .W22TO9(-4833), .W22TO10(18930), .W22TO11(3792), .W22TO12(-15472), .W22TO13(11302), .W22TO14(18666), .W22TO15(-15687), .W22TO16(7593), .W22TO17(-9782), .W22TO18(-18523), .W22TO19(-10287), .W22TO20(583), .W22TO21(-16120), .W22TO22(13946), .W22TO23(6716), .W22TO24(-6246), .W22TO25(-9470), .W22TO26(-8463), .W22TO27(11131), .W22TO28(911), .W22TO29(6716), .W22TO30(13742), .W22TO31(-10268), .W22TO32(20415), .W22TO33(10137), .W22TO34(5765), .W22TO35(3245), .W22TO36(-89), .W22TO37(11552), .W22TO38(-4412), .W22TO39(10139), .W22TO40(-13826), .W22TO41(19708), .W22TO42(1781), .W22TO43(17340), .W22TO44(-3340), .W22TO45(-4345), .W22TO46(7814), .W22TO47(14530), .W22TO48(-14715), .W22TO49(10470), .W22TO50(-6522), .W22TO51(-9747), .W22TO52(7041), .W22TO53(-9609), .W22TO54(-5415), .W22TO55(8181), .W22TO56(-12766), .W22TO57(9735), .W22TO58(-8698), .W22TO59(8997), .W22TO60(-3741), .W22TO61(22061), .W22TO62(-18829), .W22TO63(3516), .W22TO64(17471), .W22TO65(-9015), .W22TO66(-3553), .W22TO67(-9175), .W22TO68(10473), .W22TO69(19078), .W22TO70(-1704), .W22TO71(-93), .W22TO72(-10103), .W22TO73(12656), .W22TO74(-14121), .W22TO75(-6973), .W22TO76(12210), .W22TO77(-17927), .W22TO78(3959), .W22TO79(-5941), .W22TO80(-8884), .W22TO81(14758), .W22TO82(1111), .W22TO83(-13688), .W22TO84(13616), .W22TO85(-10762), .W22TO86(12075), .W22TO87(-11332), .W22TO88(-2808), .W22TO89(10517), .W22TO90(7118), .W22TO91(2387), .W22TO92(8865), .W22TO93(-9136), .W22TO94(-15226), .W22TO95(11327), .W22TO96(17901), .W22TO97(-17606), .W22TO98(-2727), .W22TO99(-900), .W23TO0(-15762), .W23TO1(10182), .W23TO2(15567), .W23TO3(-3751), .W23TO4(-18200), .W23TO5(-1309), .W23TO6(8827), .W23TO7(-6273), .W23TO8(10946), .W23TO9(-5076), .W23TO10(12508), .W23TO11(-5700), .W23TO12(-12394), .W23TO13(-5353), .W23TO14(3014), .W23TO15(-15126), .W23TO16(-14509), .W23TO17(-1916), .W23TO18(-7168), .W23TO19(-9862), .W23TO20(-2438), .W23TO21(-261), .W23TO22(2456), .W23TO23(15270), .W23TO24(-1227), .W23TO25(-2212), .W23TO26(-10114), .W23TO27(7266), .W23TO28(-18801), .W23TO29(-11970), .W23TO30(-4401), .W23TO31(15101), .W23TO32(11800), .W23TO33(-12011), .W23TO34(18557), .W23TO35(-5319), .W23TO36(-3477), .W23TO37(18550), .W23TO38(14312), .W23TO39(-12352), .W23TO40(2417), .W23TO41(-8715), .W23TO42(-14092), .W23TO43(-970), .W23TO44(-939), .W23TO45(15141), .W23TO46(14261), .W23TO47(-16908), .W23TO48(981), .W23TO49(2623), .W23TO50(-9658), .W23TO51(-12197), .W23TO52(1804), .W23TO53(17026), .W23TO54(-3926), .W23TO55(-7351), .W23TO56(6961), .W23TO57(5223), .W23TO58(-5996), .W23TO59(6531), .W23TO60(-11929), .W23TO61(4780), .W23TO62(-11792), .W23TO63(14723), .W23TO64(11192), .W23TO65(9785), .W23TO66(12341), .W23TO67(-6889), .W23TO68(12302), .W23TO69(-8233), .W23TO70(3068), .W23TO71(9304), .W23TO72(-12672), .W23TO73(-17959), .W23TO74(1851), .W23TO75(-10305), .W23TO76(15451), .W23TO77(17711), .W23TO78(-4333), .W23TO79(17439), .W23TO80(-1163), .W23TO81(-9142), .W23TO82(-3451), .W23TO83(13374), .W23TO84(675), .W23TO85(-4439), .W23TO86(6956), .W23TO87(-7352), .W23TO88(-12082), .W23TO89(11924), .W23TO90(-3519), .W23TO91(-5635), .W23TO92(18559), .W23TO93(18908), .W23TO94(7352), .W23TO95(12222), .W23TO96(6717), .W23TO97(-2154), .W23TO98(-10427), .W23TO99(565), .W24TO0(-18506), .W24TO1(514), .W24TO2(4797), .W24TO3(1012), .W24TO4(-2967), .W24TO5(-12192), .W24TO6(5461), .W24TO7(-4860), .W24TO8(10577), .W24TO9(-17937), .W24TO10(-15535), .W24TO11(14920), .W24TO12(-9488), .W24TO13(-9585), .W24TO14(-18468), .W24TO15(-2702), .W24TO16(1521), .W24TO17(1688), .W24TO18(18637), .W24TO19(-13517), .W24TO20(-14115), .W24TO21(-3091), .W24TO22(3034), .W24TO23(2006), .W24TO24(9990), .W24TO25(-3221), .W24TO26(-4064), .W24TO27(7483), .W24TO28(-18834), .W24TO29(7220), .W24TO30(8225), .W24TO31(16908), .W24TO32(7490), .W24TO33(-1678), .W24TO34(-17522), .W24TO35(787), .W24TO36(-17742), .W24TO37(16373), .W24TO38(10261), .W24TO39(-1152), .W24TO40(-11675), .W24TO41(7917), .W24TO42(-3145), .W24TO43(-5812), .W24TO44(-3229), .W24TO45(3518), .W24TO46(5166), .W24TO47(16532), .W24TO48(-14088), .W24TO49(-1764), .W24TO50(8141), .W24TO51(8007), .W24TO52(16355), .W24TO53(-4614), .W24TO54(18605), .W24TO55(-11239), .W24TO56(5647), .W24TO57(16840), .W24TO58(5309), .W24TO59(9412), .W24TO60(-6158), .W24TO61(-17987), .W24TO62(-10613), .W24TO63(-6656), .W24TO64(-11768), .W24TO65(-6368), .W24TO66(11452), .W24TO67(-6395), .W24TO68(-572), .W24TO69(14903), .W24TO70(14480), .W24TO71(-11430), .W24TO72(9941), .W24TO73(-1981), .W24TO74(2686), .W24TO75(9126), .W24TO76(4777), .W24TO77(16815), .W24TO78(11530), .W24TO79(-8200), .W24TO80(-1414), .W24TO81(-12398), .W24TO82(-7324), .W24TO83(12084), .W24TO84(-10055), .W24TO85(-18732), .W24TO86(13580), .W24TO87(-717), .W24TO88(14916), .W24TO89(18681), .W24TO90(31), .W24TO91(-4300), .W24TO92(-13175), .W24TO93(-9056), .W24TO94(-14974), .W24TO95(-9444), .W24TO96(-5647), .W24TO97(-19131), .W24TO98(613), .W24TO99(15317), .W25TO0(-16063), .W25TO1(13255), .W25TO2(-791), .W25TO3(11152), .W25TO4(-20206), .W25TO5(11646), .W25TO6(8682), .W25TO7(2388), .W25TO8(-12652), .W25TO9(-7580), .W25TO10(-2260), .W25TO11(9411), .W25TO12(14127), .W25TO13(-18997), .W25TO14(1934), .W25TO15(-4400), .W25TO16(18358), .W25TO17(3393), .W25TO18(-3265), .W25TO19(-9396), .W25TO20(17980), .W25TO21(182), .W25TO22(-8256), .W25TO23(7617), .W25TO24(-12132), .W25TO25(-2814), .W25TO26(-11080), .W25TO27(16052), .W25TO28(-15943), .W25TO29(-7812), .W25TO30(-11700), .W25TO31(9198), .W25TO32(4587), .W25TO33(1964), .W25TO34(-849), .W25TO35(-14422), .W25TO36(16015), .W25TO37(-7559), .W25TO38(9254), .W25TO39(-3166), .W25TO40(8360), .W25TO41(6816), .W25TO42(-18049), .W25TO43(-9099), .W25TO44(-10898), .W25TO45(-15186), .W25TO46(-7223), .W25TO47(-12055), .W25TO48(-16177), .W25TO49(-11727), .W25TO50(-18994), .W25TO51(12610), .W25TO52(-18832), .W25TO53(-12458), .W25TO54(-4875), .W25TO55(-5066), .W25TO56(19419), .W25TO57(440), .W25TO58(-13351), .W25TO59(7170), .W25TO60(9122), .W25TO61(2971), .W25TO62(8841), .W25TO63(-8993), .W25TO64(-2241), .W25TO65(-10243), .W25TO66(-17865), .W25TO67(-3551), .W25TO68(-6862), .W25TO69(11740), .W25TO70(8189), .W25TO71(4817), .W25TO72(6722), .W25TO73(4785), .W25TO74(-5222), .W25TO75(-29), .W25TO76(19304), .W25TO77(-19885), .W25TO78(10194), .W25TO79(-14230), .W25TO80(-800), .W25TO81(-5167), .W25TO82(-17909), .W25TO83(6499), .W25TO84(606), .W25TO85(-9083), .W25TO86(12792), .W25TO87(14779), .W25TO88(-7103), .W25TO89(-16440), .W25TO90(8231), .W25TO91(13462), .W25TO92(6371), .W25TO93(558), .W25TO94(-8195), .W25TO95(-19320), .W25TO96(5447), .W25TO97(17804), .W25TO98(9271), .W25TO99(-3902), .W26TO0(-12453), .W26TO1(-2093), .W26TO2(-12173), .W26TO3(16499), .W26TO4(3077), .W26TO5(15194), .W26TO6(11385), .W26TO7(-23719), .W26TO8(-14569), .W26TO9(15025), .W26TO10(13132), .W26TO11(14025), .W26TO12(-8949), .W26TO13(-2558), .W26TO14(15842), .W26TO15(2687), .W26TO16(15733), .W26TO17(-6723), .W26TO18(-11911), .W26TO19(-19777), .W26TO20(-5938), .W26TO21(-14350), .W26TO22(11193), .W26TO23(-15304), .W26TO24(-25968), .W26TO25(5811), .W26TO26(7180), .W26TO27(-4316), .W26TO28(-10784), .W26TO29(12840), .W26TO30(-10700), .W26TO31(4282), .W26TO32(4674), .W26TO33(-2747), .W26TO34(-4656), .W26TO35(6413), .W26TO36(-2895), .W26TO37(-5634), .W26TO38(-15304), .W26TO39(9363), .W26TO40(-5559), .W26TO41(333), .W26TO42(8608), .W26TO43(7980), .W26TO44(11562), .W26TO45(-15632), .W26TO46(-4106), .W26TO47(-8140), .W26TO48(4409), .W26TO49(19244), .W26TO50(-13474), .W26TO51(-3634), .W26TO52(8609), .W26TO53(-6951), .W26TO54(17555), .W26TO55(-19826), .W26TO56(-3825), .W26TO57(2858), .W26TO58(3646), .W26TO59(-24141), .W26TO60(14498), .W26TO61(-14380), .W26TO62(-12386), .W26TO63(6745), .W26TO64(-8546), .W26TO65(-9968), .W26TO66(-20707), .W26TO67(-9434), .W26TO68(773), .W26TO69(3205), .W26TO70(-19560), .W26TO71(11027), .W26TO72(-7072), .W26TO73(6110), .W26TO74(6288), .W26TO75(4360), .W26TO76(-14569), .W26TO77(9548), .W26TO78(8070), .W26TO79(-20495), .W26TO80(-3648), .W26TO81(17167), .W26TO82(6182), .W26TO83(-16662), .W26TO84(-10687), .W26TO85(12591), .W26TO86(6353), .W26TO87(10248), .W26TO88(7866), .W26TO89(-12717), .W26TO90(18835), .W26TO91(-29922), .W26TO92(10228), .W26TO93(-25814), .W26TO94(-10662), .W26TO95(-13665), .W26TO96(-647), .W26TO97(-3345), .W26TO98(3499), .W26TO99(-8412), .W27TO0(-6409), .W27TO1(8001), .W27TO2(-4754), .W27TO3(-5253), .W27TO4(-12557), .W27TO5(-8631), .W27TO6(9661), .W27TO7(1258), .W27TO8(22690), .W27TO9(-6585), .W27TO10(16696), .W27TO11(-14085), .W27TO12(13724), .W27TO13(12983), .W27TO14(-19074), .W27TO15(1278), .W27TO16(-7386), .W27TO17(4665), .W27TO18(-2865), .W27TO19(6584), .W27TO20(-8375), .W27TO21(13915), .W27TO22(6966), .W27TO23(-1453), .W27TO24(-4744), .W27TO25(14859), .W27TO26(-2759), .W27TO27(4282), .W27TO28(-6898), .W27TO29(-12184), .W27TO30(9435), .W27TO31(5680), .W27TO32(-11312), .W27TO33(-1426), .W27TO34(-11887), .W27TO35(6388), .W27TO36(3241), .W27TO37(4546), .W27TO38(-17718), .W27TO39(6451), .W27TO40(-4405), .W27TO41(-2467), .W27TO42(11049), .W27TO43(-4374), .W27TO44(9933), .W27TO45(-703), .W27TO46(-11226), .W27TO47(980), .W27TO48(11452), .W27TO49(15772), .W27TO50(-9134), .W27TO51(2462), .W27TO52(-16022), .W27TO53(-10095), .W27TO54(-12968), .W27TO55(15241), .W27TO56(966), .W27TO57(-6000), .W27TO58(-22644), .W27TO59(-27394), .W27TO60(-3056), .W27TO61(-7595), .W27TO62(13229), .W27TO63(17268), .W27TO64(-7246), .W27TO65(-4701), .W27TO66(5584), .W27TO67(2568), .W27TO68(16461), .W27TO69(-6465), .W27TO70(11817), .W27TO71(17573), .W27TO72(-12982), .W27TO73(3441), .W27TO74(16543), .W27TO75(-14608), .W27TO76(-6930), .W27TO77(-13563), .W27TO78(-27180), .W27TO79(-2671), .W27TO80(3139), .W27TO81(-3209), .W27TO82(16661), .W27TO83(2237), .W27TO84(22271), .W27TO85(10880), .W27TO86(2880), .W27TO87(17621), .W27TO88(18261), .W27TO89(-11967), .W27TO90(-3858), .W27TO91(-4702), .W27TO92(-12611), .W27TO93(-3594), .W27TO94(-318), .W27TO95(-10456), .W27TO96(10622), .W27TO97(-7987), .W27TO98(-15425), .W27TO99(-5428), .W28TO0(-4805), .W28TO1(-5805), .W28TO2(-28356), .W28TO3(-20582), .W28TO4(-21114), .W28TO5(3614), .W28TO6(-601), .W28TO7(4575), .W28TO8(-11398), .W28TO9(-371), .W28TO10(-16670), .W28TO11(9528), .W28TO12(15077), .W28TO13(7211), .W28TO14(-8180), .W28TO15(5575), .W28TO16(14695), .W28TO17(3007), .W28TO18(21677), .W28TO19(-14422), .W28TO20(13167), .W28TO21(-16848), .W28TO22(-9192), .W28TO23(13980), .W28TO24(-12997), .W28TO25(9680), .W28TO26(-9720), .W28TO27(-10626), .W28TO28(4431), .W28TO29(13322), .W28TO30(-4329), .W28TO31(-2572), .W28TO32(1093), .W28TO33(-11862), .W28TO34(2303), .W28TO35(9348), .W28TO36(3962), .W28TO37(7861), .W28TO38(-12994), .W28TO39(-11357), .W28TO40(3264), .W28TO41(-15165), .W28TO42(6981), .W28TO43(-14988), .W28TO44(7912), .W28TO45(4671), .W28TO46(-12736), .W28TO47(7257), .W28TO48(13456), .W28TO49(10055), .W28TO50(3656), .W28TO51(-15016), .W28TO52(-8031), .W28TO53(16592), .W28TO54(-12589), .W28TO55(-8209), .W28TO56(15302), .W28TO57(10449), .W28TO58(6576), .W28TO59(-6589), .W28TO60(-1874), .W28TO61(9898), .W28TO62(4090), .W28TO63(-2628), .W28TO64(3791), .W28TO65(4034), .W28TO66(-4892), .W28TO67(-4342), .W28TO68(9355), .W28TO69(84), .W28TO70(-2878), .W28TO71(10119), .W28TO72(-10288), .W28TO73(-20547), .W28TO74(1500), .W28TO75(-11567), .W28TO76(-8706), .W28TO77(-2635), .W28TO78(-9671), .W28TO79(6827), .W28TO80(-16527), .W28TO81(16093), .W28TO82(25237), .W28TO83(3639), .W28TO84(181), .W28TO85(-4844), .W28TO86(-8594), .W28TO87(2656), .W28TO88(4105), .W28TO89(8775), .W28TO90(7967), .W28TO91(-4038), .W28TO92(16173), .W28TO93(5457), .W28TO94(-3299), .W28TO95(26328), .W28TO96(-10828), .W28TO97(3370), .W28TO98(7708), .W28TO99(-6002), .W29TO0(-12031), .W29TO1(-5836), .W29TO2(19483), .W29TO3(-5418), .W29TO4(-11894), .W29TO5(-6486), .W29TO6(14750), .W29TO7(1923), .W29TO8(-5934), .W29TO9(5340), .W29TO10(13245), .W29TO11(-551), .W29TO12(-34), .W29TO13(17219), .W29TO14(-16173), .W29TO15(17658), .W29TO16(25502), .W29TO17(-5814), .W29TO18(-2461), .W29TO19(-1703), .W29TO20(3149), .W29TO21(5802), .W29TO22(16417), .W29TO23(-13388), .W29TO24(-13472), .W29TO25(2423), .W29TO26(2541), .W29TO27(-16891), .W29TO28(-2732), .W29TO29(17301), .W29TO30(-4695), .W29TO31(-12414), .W29TO32(7082), .W29TO33(-166), .W29TO34(-8168), .W29TO35(-1581), .W29TO36(-13611), .W29TO37(4029), .W29TO38(9438), .W29TO39(8801), .W29TO40(1604), .W29TO41(-12924), .W29TO42(16038), .W29TO43(-1138), .W29TO44(-4075), .W29TO45(-18588), .W29TO46(-595), .W29TO47(9249), .W29TO48(13973), .W29TO49(11574), .W29TO50(3860), .W29TO51(12844), .W29TO52(12310), .W29TO53(-12307), .W29TO54(438), .W29TO55(-4215), .W29TO56(6913), .W29TO57(-13380), .W29TO58(-3912), .W29TO59(-11948), .W29TO60(-5557), .W29TO61(-9669), .W29TO62(-11127), .W29TO63(-6400), .W29TO64(-13231), .W29TO65(15377), .W29TO66(7097), .W29TO67(-22043), .W29TO68(-3528), .W29TO69(-7414), .W29TO70(-518), .W29TO71(-6997), .W29TO72(17054), .W29TO73(-2562), .W29TO74(3113), .W29TO75(-2172), .W29TO76(-23709), .W29TO77(5796), .W29TO78(7373), .W29TO79(-12678), .W29TO80(3366), .W29TO81(-7627), .W29TO82(-23831), .W29TO83(-2914), .W29TO84(20999), .W29TO85(20943), .W29TO86(-1930), .W29TO87(-9029), .W29TO88(-10110), .W29TO89(-12605), .W29TO90(-6572), .W29TO91(-13324), .W29TO92(20140), .W29TO93(-4156), .W29TO94(-21460), .W29TO95(-20389), .W29TO96(-13612), .W29TO97(-16251), .W29TO98(9680), .W29TO99(17035), .W30TO0(-2535), .W30TO1(-6849), .W30TO2(9229), .W30TO3(7745), .W30TO4(12319), .W30TO5(37), .W30TO6(6408), .W30TO7(-6093), .W30TO8(-3250), .W30TO9(18299), .W30TO10(-14437), .W30TO11(-10878), .W30TO12(7658), .W30TO13(-10079), .W30TO14(19149), .W30TO15(-17202), .W30TO16(9113), .W30TO17(14041), .W30TO18(6628), .W30TO19(-17924), .W30TO20(-17401), .W30TO21(-3687), .W30TO22(1076), .W30TO23(12442), .W30TO24(10267), .W30TO25(-16311), .W30TO26(-5928), .W30TO27(4880), .W30TO28(-8955), .W30TO29(24990), .W30TO30(-391), .W30TO31(14359), .W30TO32(1893), .W30TO33(-9531), .W30TO34(4788), .W30TO35(2811), .W30TO36(1445), .W30TO37(-3162), .W30TO38(8599), .W30TO39(-7181), .W30TO40(-18209), .W30TO41(2186), .W30TO42(2065), .W30TO43(-10359), .W30TO44(12355), .W30TO45(11526), .W30TO46(-18648), .W30TO47(-14403), .W30TO48(16456), .W30TO49(10151), .W30TO50(13356), .W30TO51(16335), .W30TO52(-9098), .W30TO53(-6550), .W30TO54(18853), .W30TO55(-3449), .W30TO56(-1933), .W30TO57(2515), .W30TO58(-1109), .W30TO59(-18421), .W30TO60(4432), .W30TO61(3216), .W30TO62(15632), .W30TO63(-13035), .W30TO64(5535), .W30TO65(6276), .W30TO66(-8476), .W30TO67(-11232), .W30TO68(11804), .W30TO69(3924), .W30TO70(9958), .W30TO71(11536), .W30TO72(5666), .W30TO73(-9431), .W30TO74(-8270), .W30TO75(12855), .W30TO76(-763), .W30TO77(14573), .W30TO78(21272), .W30TO79(-1711), .W30TO80(8807), .W30TO81(-885), .W30TO82(-22008), .W30TO83(8679), .W30TO84(6309), .W30TO85(16560), .W30TO86(13575), .W30TO87(13751), .W30TO88(-7443), .W30TO89(-9021), .W30TO90(16878), .W30TO91(-5233), .W30TO92(19007), .W30TO93(-5792), .W30TO94(10056), .W30TO95(414), .W30TO96(1366), .W30TO97(-13340), .W30TO98(15051), .W30TO99(-18003), .W31TO0(-6529), .W31TO1(-10609), .W31TO2(-15534), .W31TO3(5948), .W31TO4(14147), .W31TO5(-5921), .W31TO6(-2298), .W31TO7(7288), .W31TO8(-7061), .W31TO9(-15785), .W31TO10(1441), .W31TO11(15653), .W31TO12(87), .W31TO13(10419), .W31TO14(5426), .W31TO15(-2174), .W31TO16(452), .W31TO17(-15545), .W31TO18(-17469), .W31TO19(-11969), .W31TO20(-17847), .W31TO21(-7069), .W31TO22(-5594), .W31TO23(-14911), .W31TO24(5607), .W31TO25(8031), .W31TO26(-3112), .W31TO27(-10176), .W31TO28(-1535), .W31TO29(-6052), .W31TO30(-2974), .W31TO31(7787), .W31TO32(1553), .W31TO33(8879), .W31TO34(-16391), .W31TO35(8846), .W31TO36(10617), .W31TO37(14683), .W31TO38(14930), .W31TO39(5301), .W31TO40(-6821), .W31TO41(5672), .W31TO42(-11356), .W31TO43(9110), .W31TO44(3539), .W31TO45(4369), .W31TO46(-12341), .W31TO47(-2782), .W31TO48(-9668), .W31TO49(-8338), .W31TO50(18486), .W31TO51(46), .W31TO52(-15496), .W31TO53(-15212), .W31TO54(14832), .W31TO55(-12503), .W31TO56(352), .W31TO57(4084), .W31TO58(-18955), .W31TO59(-8984), .W31TO60(-13747), .W31TO61(-9733), .W31TO62(-18119), .W31TO63(14898), .W31TO64(9875), .W31TO65(4200), .W31TO66(16147), .W31TO67(14023), .W31TO68(-4029), .W31TO69(10250), .W31TO70(12542), .W31TO71(17666), .W31TO72(3707), .W31TO73(-3309), .W31TO74(11107), .W31TO75(-17652), .W31TO76(-9644), .W31TO77(2826), .W31TO78(-17355), .W31TO79(15458), .W31TO80(-15137), .W31TO81(16563), .W31TO82(18671), .W31TO83(-11739), .W31TO84(-4089), .W31TO85(9124), .W31TO86(15703), .W31TO87(16905), .W31TO88(-18534), .W31TO89(-10747), .W31TO90(8719), .W31TO91(366), .W31TO92(11387), .W31TO93(-7253), .W31TO94(11688), .W31TO95(8438), .W31TO96(-7778), .W31TO97(-18741), .W31TO98(-7744), .W31TO99(-6304), .W32TO0(9061), .W32TO1(-11255), .W32TO2(-11200), .W32TO3(-5964), .W32TO4(-14558), .W32TO5(12724), .W32TO6(-17891), .W32TO7(-18938), .W32TO8(-6463), .W32TO9(-7994), .W32TO10(18638), .W32TO11(27), .W32TO12(-3969), .W32TO13(14142), .W32TO14(5986), .W32TO15(-249), .W32TO16(-16795), .W32TO17(1483), .W32TO18(9282), .W32TO19(13818), .W32TO20(-10917), .W32TO21(5011), .W32TO22(16857), .W32TO23(10264), .W32TO24(10724), .W32TO25(-480), .W32TO26(-351), .W32TO27(-12033), .W32TO28(3451), .W32TO29(-6565), .W32TO30(2794), .W32TO31(-6996), .W32TO32(-18874), .W32TO33(10890), .W32TO34(-6170), .W32TO35(-11675), .W32TO36(15748), .W32TO37(-9383), .W32TO38(-17633), .W32TO39(16273), .W32TO40(-15848), .W32TO41(-5874), .W32TO42(9908), .W32TO43(-14024), .W32TO44(-17207), .W32TO45(-10227), .W32TO46(-4100), .W32TO47(-14927), .W32TO48(-4395), .W32TO49(-5053), .W32TO50(15497), .W32TO51(-1501), .W32TO52(-1018), .W32TO53(15976), .W32TO54(-15117), .W32TO55(-13625), .W32TO56(15807), .W32TO57(-10526), .W32TO58(-17228), .W32TO59(-6462), .W32TO60(7516), .W32TO61(-12443), .W32TO62(-17753), .W32TO63(7705), .W32TO64(-10366), .W32TO65(-812), .W32TO66(15618), .W32TO67(-11143), .W32TO68(-11837), .W32TO69(12573), .W32TO70(11088), .W32TO71(-14195), .W32TO72(-18628), .W32TO73(9534), .W32TO74(-8069), .W32TO75(-6271), .W32TO76(9649), .W32TO77(7274), .W32TO78(10249), .W32TO79(-12960), .W32TO80(-3811), .W32TO81(3753), .W32TO82(1902), .W32TO83(18689), .W32TO84(-2697), .W32TO85(2711), .W32TO86(10571), .W32TO87(7242), .W32TO88(-12173), .W32TO89(3586), .W32TO90(-16480), .W32TO91(14450), .W32TO92(-3782), .W32TO93(-10256), .W32TO94(10071), .W32TO95(17963), .W32TO96(-8295), .W32TO97(-2400), .W32TO98(-13815), .W32TO99(1106), .W33TO0(17426), .W33TO1(-12656), .W33TO2(11440), .W33TO3(-3256), .W33TO4(-4998), .W33TO5(-13420), .W33TO6(-12415), .W33TO7(-13072), .W33TO8(10477), .W33TO9(5801), .W33TO10(17131), .W33TO11(-12061), .W33TO12(7674), .W33TO13(-21071), .W33TO14(-14538), .W33TO15(5970), .W33TO16(-5918), .W33TO17(16314), .W33TO18(-13506), .W33TO19(-12023), .W33TO20(-15122), .W33TO21(-1912), .W33TO22(-22230), .W33TO23(608), .W33TO24(-13918), .W33TO25(-6825), .W33TO26(-8452), .W33TO27(-18138), .W33TO28(-155), .W33TO29(11249), .W33TO30(-13201), .W33TO31(-8455), .W33TO32(-15645), .W33TO33(2889), .W33TO34(11546), .W33TO35(-6390), .W33TO36(-7513), .W33TO37(1647), .W33TO38(18025), .W33TO39(1984), .W33TO40(2481), .W33TO41(1401), .W33TO42(5483), .W33TO43(-13324), .W33TO44(-18388), .W33TO45(-201), .W33TO46(-13765), .W33TO47(-19605), .W33TO48(11192), .W33TO49(13569), .W33TO50(2618), .W33TO51(-13945), .W33TO52(1702), .W33TO53(-10434), .W33TO54(5429), .W33TO55(3020), .W33TO56(17779), .W33TO57(7619), .W33TO58(-9265), .W33TO59(12478), .W33TO60(8657), .W33TO61(9585), .W33TO62(-6041), .W33TO63(-18427), .W33TO64(-6430), .W33TO65(-6388), .W33TO66(-13388), .W33TO67(-11891), .W33TO68(-8327), .W33TO69(10052), .W33TO70(-20497), .W33TO71(-7498), .W33TO72(-9921), .W33TO73(-11042), .W33TO74(-378), .W33TO75(17387), .W33TO76(7917), .W33TO77(-16278), .W33TO78(612), .W33TO79(-16433), .W33TO80(-7138), .W33TO81(-4946), .W33TO82(-27368), .W33TO83(-19945), .W33TO84(-615), .W33TO85(9969), .W33TO86(-5809), .W33TO87(17222), .W33TO88(-4100), .W33TO89(9314), .W33TO90(-17319), .W33TO91(10358), .W33TO92(-9603), .W33TO93(6431), .W33TO94(-20010), .W33TO95(-8969), .W33TO96(2515), .W33TO97(-14353), .W33TO98(-3106), .W33TO99(-18014), .W34TO0(-6012), .W34TO1(-3092), .W34TO2(-16363), .W34TO3(-18256), .W34TO4(9207), .W34TO5(-10566), .W34TO6(-15723), .W34TO7(-964), .W34TO8(21698), .W34TO9(11686), .W34TO10(9570), .W34TO11(1405), .W34TO12(2785), .W34TO13(-10868), .W34TO14(-18330), .W34TO15(-1178), .W34TO16(9400), .W34TO17(-15331), .W34TO18(3380), .W34TO19(-12445), .W34TO20(-5007), .W34TO21(-14387), .W34TO22(-22609), .W34TO23(8064), .W34TO24(-22207), .W34TO25(-21074), .W34TO26(13209), .W34TO27(3701), .W34TO28(6687), .W34TO29(2139), .W34TO30(1751), .W34TO31(15008), .W34TO32(-4933), .W34TO33(11904), .W34TO34(-18982), .W34TO35(13000), .W34TO36(-8835), .W34TO37(9790), .W34TO38(10382), .W34TO39(18305), .W34TO40(-2228), .W34TO41(-4545), .W34TO42(10817), .W34TO43(7038), .W34TO44(15717), .W34TO45(11227), .W34TO46(13470), .W34TO47(4900), .W34TO48(5457), .W34TO49(-5640), .W34TO50(11244), .W34TO51(6981), .W34TO52(4140), .W34TO53(-2136), .W34TO54(3322), .W34TO55(-6390), .W34TO56(1618), .W34TO57(-14367), .W34TO58(-4547), .W34TO59(-4481), .W34TO60(5146), .W34TO61(-952), .W34TO62(12755), .W34TO63(17438), .W34TO64(-8976), .W34TO65(11312), .W34TO66(8175), .W34TO67(3222), .W34TO68(-9549), .W34TO69(17917), .W34TO70(-6196), .W34TO71(5148), .W34TO72(11857), .W34TO73(2815), .W34TO74(6849), .W34TO75(-14307), .W34TO76(12595), .W34TO77(16790), .W34TO78(10250), .W34TO79(-15465), .W34TO80(-9199), .W34TO81(15774), .W34TO82(3531), .W34TO83(-12149), .W34TO84(-2845), .W34TO85(12413), .W34TO86(10699), .W34TO87(-1093), .W34TO88(6990), .W34TO89(-192), .W34TO90(13198), .W34TO91(-196), .W34TO92(-14604), .W34TO93(-8349), .W34TO94(11330), .W34TO95(12212), .W34TO96(4325), .W34TO97(12709), .W34TO98(-4906), .W34TO99(9976), .W35TO0(5172), .W35TO1(-1257), .W35TO2(-11217), .W35TO3(15485), .W35TO4(-14688), .W35TO5(11764), .W35TO6(-3337), .W35TO7(14306), .W35TO8(18913), .W35TO9(12827), .W35TO10(2915), .W35TO11(7215), .W35TO12(-18066), .W35TO13(-3496), .W35TO14(15018), .W35TO15(13943), .W35TO16(1833), .W35TO17(5659), .W35TO18(-8790), .W35TO19(-640), .W35TO20(-19217), .W35TO21(-16920), .W35TO22(-7713), .W35TO23(-18674), .W35TO24(13310), .W35TO25(-16384), .W35TO26(7430), .W35TO27(313), .W35TO28(4770), .W35TO29(11862), .W35TO30(6398), .W35TO31(15880), .W35TO32(12867), .W35TO33(15692), .W35TO34(-19406), .W35TO35(-1766), .W35TO36(16551), .W35TO37(-874), .W35TO38(17538), .W35TO39(-8934), .W35TO40(-21115), .W35TO41(5818), .W35TO42(-9192), .W35TO43(8721), .W35TO44(-16092), .W35TO45(-3606), .W35TO46(2360), .W35TO47(8035), .W35TO48(-20932), .W35TO49(13095), .W35TO50(22050), .W35TO51(17810), .W35TO52(-1279), .W35TO53(22912), .W35TO54(8499), .W35TO55(22179), .W35TO56(20244), .W35TO57(7729), .W35TO58(-8730), .W35TO59(1885), .W35TO60(15139), .W35TO61(1743), .W35TO62(12229), .W35TO63(-8670), .W35TO64(-186), .W35TO65(-2573), .W35TO66(-8330), .W35TO67(-17450), .W35TO68(11777), .W35TO69(19966), .W35TO70(12627), .W35TO71(-1728), .W35TO72(-6903), .W35TO73(-18465), .W35TO74(10572), .W35TO75(3051), .W35TO76(3635), .W35TO77(-10417), .W35TO78(-18985), .W35TO79(8459), .W35TO80(-463), .W35TO81(-8778), .W35TO82(-409), .W35TO83(3734), .W35TO84(3312), .W35TO85(14574), .W35TO86(-14384), .W35TO87(-553), .W35TO88(16594), .W35TO89(8430), .W35TO90(-7517), .W35TO91(2389), .W35TO92(-4773), .W35TO93(21069), .W35TO94(3669), .W35TO95(-5947), .W35TO96(-4123), .W35TO97(-14327), .W35TO98(7535), .W35TO99(6409), .W36TO0(6798), .W36TO1(4197), .W36TO2(-17393), .W36TO3(-7829), .W36TO4(-10746), .W36TO5(-9148), .W36TO6(-8094), .W36TO7(5122), .W36TO8(14509), .W36TO9(-6262), .W36TO10(2965), .W36TO11(693), .W36TO12(-9071), .W36TO13(-9063), .W36TO14(-15302), .W36TO15(-6475), .W36TO16(12005), .W36TO17(10711), .W36TO18(12507), .W36TO19(11531), .W36TO20(1863), .W36TO21(1370), .W36TO22(-9490), .W36TO23(-9722), .W36TO24(10908), .W36TO25(16086), .W36TO26(-8680), .W36TO27(5744), .W36TO28(16409), .W36TO29(-12300), .W36TO30(14668), .W36TO31(10640), .W36TO32(-5125), .W36TO33(7381), .W36TO34(-9758), .W36TO35(13679), .W36TO36(2662), .W36TO37(4391), .W36TO38(11130), .W36TO39(2149), .W36TO40(-16112), .W36TO41(7061), .W36TO42(-15360), .W36TO43(-4078), .W36TO44(5630), .W36TO45(14472), .W36TO46(-14689), .W36TO47(1088), .W36TO48(2260), .W36TO49(-13397), .W36TO50(5961), .W36TO51(3115), .W36TO52(-18129), .W36TO53(1180), .W36TO54(-10700), .W36TO55(-548), .W36TO56(-11510), .W36TO57(-2008), .W36TO58(877), .W36TO59(-9114), .W36TO60(1959), .W36TO61(-1484), .W36TO62(-12873), .W36TO63(-13880), .W36TO64(394), .W36TO65(4215), .W36TO66(-21494), .W36TO67(-1329), .W36TO68(-10989), .W36TO69(-14165), .W36TO70(8968), .W36TO71(-2129), .W36TO72(-3924), .W36TO73(12377), .W36TO74(-2980), .W36TO75(-12642), .W36TO76(359), .W36TO77(17513), .W36TO78(13985), .W36TO79(16896), .W36TO80(-10506), .W36TO81(-507), .W36TO82(-3131), .W36TO83(-20400), .W36TO84(-1925), .W36TO85(1035), .W36TO86(14792), .W36TO87(-8292), .W36TO88(13952), .W36TO89(-15680), .W36TO90(17742), .W36TO91(21272), .W36TO92(-1860), .W36TO93(20068), .W36TO94(-10120), .W36TO95(13186), .W36TO96(4991), .W36TO97(-10953), .W36TO98(-12360), .W36TO99(-4480), .W37TO0(-15672), .W37TO1(13834), .W37TO2(-19102), .W37TO3(-14340), .W37TO4(-4578), .W37TO5(11511), .W37TO6(15101), .W37TO7(-6524), .W37TO8(-6643), .W37TO9(13444), .W37TO10(18004), .W37TO11(-18210), .W37TO12(2426), .W37TO13(-9489), .W37TO14(15863), .W37TO15(16038), .W37TO16(20524), .W37TO17(-4841), .W37TO18(-4621), .W37TO19(2132), .W37TO20(2831), .W37TO21(8517), .W37TO22(11146), .W37TO23(-14069), .W37TO24(-13868), .W37TO25(12817), .W37TO26(14799), .W37TO27(-13205), .W37TO28(8397), .W37TO29(400), .W37TO30(-1614), .W37TO31(1261), .W37TO32(19253), .W37TO33(4163), .W37TO34(-18971), .W37TO35(10516), .W37TO36(-20145), .W37TO37(2842), .W37TO38(-6055), .W37TO39(6401), .W37TO40(-23133), .W37TO41(-10615), .W37TO42(756), .W37TO43(4362), .W37TO44(6290), .W37TO45(11288), .W37TO46(-14594), .W37TO47(-7145), .W37TO48(-5370), .W37TO49(-7072), .W37TO50(14049), .W37TO51(21859), .W37TO52(-557), .W37TO53(2862), .W37TO54(27399), .W37TO55(12013), .W37TO56(5845), .W37TO57(-9721), .W37TO58(-16199), .W37TO59(3340), .W37TO60(9406), .W37TO61(-11994), .W37TO62(-18323), .W37TO63(8965), .W37TO64(-17795), .W37TO65(-5099), .W37TO66(9917), .W37TO67(5274), .W37TO68(14417), .W37TO69(-15568), .W37TO70(-16173), .W37TO71(-4331), .W37TO72(-2293), .W37TO73(-10274), .W37TO74(-13175), .W37TO75(-9924), .W37TO76(-9374), .W37TO77(7754), .W37TO78(-335), .W37TO79(7149), .W37TO80(-16358), .W37TO81(10017), .W37TO82(-14719), .W37TO83(5243), .W37TO84(14099), .W37TO85(-10728), .W37TO86(7457), .W37TO87(-10049), .W37TO88(1044), .W37TO89(-8237), .W37TO90(11483), .W37TO91(20629), .W37TO92(-1911), .W37TO93(847), .W37TO94(-17121), .W37TO95(15754), .W37TO96(1221), .W37TO97(-3557), .W37TO98(-7087), .W37TO99(12413), .W38TO0(-14838), .W38TO1(-5159), .W38TO2(-5514), .W38TO3(-7514), .W38TO4(-7946), .W38TO5(3246), .W38TO6(-18223), .W38TO7(5622), .W38TO8(6928), .W38TO9(12502), .W38TO10(-11194), .W38TO11(-11669), .W38TO12(11464), .W38TO13(4139), .W38TO14(2178), .W38TO15(15809), .W38TO16(-899), .W38TO17(95), .W38TO18(15805), .W38TO19(2074), .W38TO20(-2097), .W38TO21(-5897), .W38TO22(-3797), .W38TO23(-17602), .W38TO24(7544), .W38TO25(10007), .W38TO26(14859), .W38TO27(-9558), .W38TO28(-12277), .W38TO29(16400), .W38TO30(-18000), .W38TO31(-8516), .W38TO32(13405), .W38TO33(8499), .W38TO34(-7768), .W38TO35(-1648), .W38TO36(6368), .W38TO37(13554), .W38TO38(-5355), .W38TO39(-1383), .W38TO40(10612), .W38TO41(-4615), .W38TO42(3792), .W38TO43(-8383), .W38TO44(18377), .W38TO45(5483), .W38TO46(5953), .W38TO47(-9097), .W38TO48(-6576), .W38TO49(-9778), .W38TO50(-11828), .W38TO51(11752), .W38TO52(4612), .W38TO53(-29636), .W38TO54(22561), .W38TO55(-5400), .W38TO56(-16753), .W38TO57(-5347), .W38TO58(-9456), .W38TO59(19700), .W38TO60(10309), .W38TO61(2086), .W38TO62(6305), .W38TO63(-7702), .W38TO64(-17462), .W38TO65(4719), .W38TO66(5892), .W38TO67(-15214), .W38TO68(-4733), .W38TO69(-12641), .W38TO70(3173), .W38TO71(20525), .W38TO72(-16081), .W38TO73(1415), .W38TO74(-16931), .W38TO75(-929), .W38TO76(61), .W38TO77(13657), .W38TO78(-7633), .W38TO79(-1987), .W38TO80(-14376), .W38TO81(18804), .W38TO82(-6335), .W38TO83(4024), .W38TO84(-3294), .W38TO85(-14501), .W38TO86(-8657), .W38TO87(321), .W38TO88(282), .W38TO89(12855), .W38TO90(-2751), .W38TO91(4962), .W38TO92(9534), .W38TO93(-5015), .W38TO94(-4901), .W38TO95(3646), .W38TO96(-10823), .W38TO97(-7526), .W38TO98(-12140), .W38TO99(15316), .W39TO0(-8645), .W39TO1(11816), .W39TO2(6425), .W39TO3(-1222), .W39TO4(858), .W39TO5(-17006), .W39TO6(13738), .W39TO7(-6423), .W39TO8(470), .W39TO9(6834), .W39TO10(-5514), .W39TO11(-18018), .W39TO12(-8734), .W39TO13(-6034), .W39TO14(2587), .W39TO15(-12827), .W39TO16(-2555), .W39TO17(-11579), .W39TO18(-8034), .W39TO19(6471), .W39TO20(13805), .W39TO21(-8343), .W39TO22(-17594), .W39TO23(7128), .W39TO24(-16152), .W39TO25(-11644), .W39TO26(-1729), .W39TO27(6592), .W39TO28(-11900), .W39TO29(-10817), .W39TO30(-17525), .W39TO31(14381), .W39TO32(12501), .W39TO33(16764), .W39TO34(-15426), .W39TO35(-9622), .W39TO36(-231), .W39TO37(-8224), .W39TO38(-6784), .W39TO39(16803), .W39TO40(-14923), .W39TO41(-10889), .W39TO42(-12175), .W39TO43(-3592), .W39TO44(-6538), .W39TO45(5994), .W39TO46(-6499), .W39TO47(-5460), .W39TO48(8657), .W39TO49(-6881), .W39TO50(13462), .W39TO51(4888), .W39TO52(14250), .W39TO53(-14085), .W39TO54(8921), .W39TO55(18400), .W39TO56(-3068), .W39TO57(2102), .W39TO58(-3955), .W39TO59(5805), .W39TO60(178), .W39TO61(-15917), .W39TO62(-10627), .W39TO63(17939), .W39TO64(-3543), .W39TO65(14999), .W39TO66(405), .W39TO67(-9396), .W39TO68(1635), .W39TO69(15412), .W39TO70(-18051), .W39TO71(-6858), .W39TO72(-10441), .W39TO73(-6350), .W39TO74(10258), .W39TO75(-3662), .W39TO76(7587), .W39TO77(16322), .W39TO78(-12715), .W39TO79(16943), .W39TO80(-18081), .W39TO81(-7366), .W39TO82(17787), .W39TO83(7472), .W39TO84(-2319), .W39TO85(-6572), .W39TO86(-18071), .W39TO87(18700), .W39TO88(-11287), .W39TO89(-9626), .W39TO90(-7060), .W39TO91(6505), .W39TO92(6673), .W39TO93(17465), .W39TO94(10143), .W39TO95(-7555), .W39TO96(9362), .W39TO97(-7274), .W39TO98(8127), .W39TO99(19029), .W40TO0(2542), .W40TO1(-2446), .W40TO2(-16210), .W40TO3(-18456), .W40TO4(10729), .W40TO5(13904), .W40TO6(7087), .W40TO7(-13485), .W40TO8(938), .W40TO9(-19010), .W40TO10(4265), .W40TO11(-15101), .W40TO12(-3219), .W40TO13(-12169), .W40TO14(11243), .W40TO15(-3988), .W40TO16(-6571), .W40TO17(14419), .W40TO18(17372), .W40TO19(6364), .W40TO20(9851), .W40TO21(-364), .W40TO22(-664), .W40TO23(2894), .W40TO24(5325), .W40TO25(11426), .W40TO26(-7318), .W40TO27(-6603), .W40TO28(13532), .W40TO29(527), .W40TO30(11805), .W40TO31(-14122), .W40TO32(4680), .W40TO33(16599), .W40TO34(5023), .W40TO35(14946), .W40TO36(-9978), .W40TO37(17905), .W40TO38(16870), .W40TO39(3140), .W40TO40(-1887), .W40TO41(-606), .W40TO42(-17197), .W40TO43(18063), .W40TO44(2655), .W40TO45(11982), .W40TO46(-15909), .W40TO47(-5197), .W40TO48(-6099), .W40TO49(-2261), .W40TO50(-1209), .W40TO51(-8270), .W40TO52(-14847), .W40TO53(-11390), .W40TO54(-17890), .W40TO55(-6928), .W40TO56(-1766), .W40TO57(2756), .W40TO58(-18887), .W40TO59(-3228), .W40TO60(10721), .W40TO61(12823), .W40TO62(7637), .W40TO63(17591), .W40TO64(-13393), .W40TO65(-13473), .W40TO66(-4120), .W40TO67(10736), .W40TO68(8179), .W40TO69(-102), .W40TO70(6303), .W40TO71(7766), .W40TO72(18623), .W40TO73(12741), .W40TO74(684), .W40TO75(-9681), .W40TO76(5132), .W40TO77(16596), .W40TO78(-3766), .W40TO79(-2522), .W40TO80(18814), .W40TO81(-18186), .W40TO82(-14430), .W40TO83(14677), .W40TO84(-621), .W40TO85(6008), .W40TO86(-15575), .W40TO87(9803), .W40TO88(9900), .W40TO89(-12016), .W40TO90(-913), .W40TO91(10519), .W40TO92(7139), .W40TO93(-18244), .W40TO94(6592), .W40TO95(5325), .W40TO96(-12594), .W40TO97(-2007), .W40TO98(13346), .W40TO99(-3920), .W41TO0(12446), .W41TO1(-5822), .W41TO2(11651), .W41TO3(14206), .W41TO4(-6425), .W41TO5(4532), .W41TO6(-15768), .W41TO7(6945), .W41TO8(-12836), .W41TO9(14694), .W41TO10(-6766), .W41TO11(-10760), .W41TO12(-10358), .W41TO13(-6146), .W41TO14(5700), .W41TO15(15998), .W41TO16(-13037), .W41TO17(-17629), .W41TO18(11646), .W41TO19(-17047), .W41TO20(-7945), .W41TO21(-14157), .W41TO22(15951), .W41TO23(7796), .W41TO24(705), .W41TO25(8436), .W41TO26(-9361), .W41TO27(-10864), .W41TO28(11193), .W41TO29(13749), .W41TO30(-19515), .W41TO31(11074), .W41TO32(-14754), .W41TO33(-19826), .W41TO34(-18926), .W41TO35(-14384), .W41TO36(16209), .W41TO37(-14124), .W41TO38(3051), .W41TO39(11278), .W41TO40(1973), .W41TO41(13276), .W41TO42(-18106), .W41TO43(7048), .W41TO44(13365), .W41TO45(10634), .W41TO46(11452), .W41TO47(-12629), .W41TO48(8886), .W41TO49(-6031), .W41TO50(18173), .W41TO51(20813), .W41TO52(-905), .W41TO53(7606), .W41TO54(1612), .W41TO55(14919), .W41TO56(329), .W41TO57(-17816), .W41TO58(-14634), .W41TO59(13647), .W41TO60(-5979), .W41TO61(-21346), .W41TO62(2512), .W41TO63(-22020), .W41TO64(-18020), .W41TO65(-12215), .W41TO66(947), .W41TO67(-9480), .W41TO68(-255), .W41TO69(-2146), .W41TO70(-17873), .W41TO71(-11378), .W41TO72(18895), .W41TO73(9181), .W41TO74(-5266), .W41TO75(3692), .W41TO76(7113), .W41TO77(-3851), .W41TO78(10098), .W41TO79(2196), .W41TO80(-194), .W41TO81(-18783), .W41TO82(-1844), .W41TO83(-973), .W41TO84(-9143), .W41TO85(-1505), .W41TO86(-2905), .W41TO87(-1018), .W41TO88(4367), .W41TO89(-17661), .W41TO90(-17176), .W41TO91(-2377), .W41TO92(2357), .W41TO93(14291), .W41TO94(5467), .W41TO95(-859), .W41TO96(-9099), .W41TO97(10964), .W41TO98(2770), .W41TO99(-3019), .W42TO0(-11859), .W42TO1(137), .W42TO2(12627), .W42TO3(15476), .W42TO4(20043), .W42TO5(-19862), .W42TO6(17361), .W42TO7(-17351), .W42TO8(-1235), .W42TO9(14651), .W42TO10(16463), .W42TO11(12782), .W42TO12(-7230), .W42TO13(752), .W42TO14(6864), .W42TO15(16346), .W42TO16(12186), .W42TO17(-17641), .W42TO18(-11085), .W42TO19(-4944), .W42TO20(-351), .W42TO21(-5552), .W42TO22(874), .W42TO23(9140), .W42TO24(-3504), .W42TO25(7884), .W42TO26(-5421), .W42TO27(-844), .W42TO28(-17506), .W42TO29(-1672), .W42TO30(14952), .W42TO31(12176), .W42TO32(-5486), .W42TO33(14052), .W42TO34(-15019), .W42TO35(-12773), .W42TO36(2026), .W42TO37(247), .W42TO38(12517), .W42TO39(2282), .W42TO40(12276), .W42TO41(28840), .W42TO42(4432), .W42TO43(9178), .W42TO44(-9813), .W42TO45(-13667), .W42TO46(-1996), .W42TO47(-10060), .W42TO48(-17287), .W42TO49(-9769), .W42TO50(10234), .W42TO51(-5486), .W42TO52(14009), .W42TO53(5877), .W42TO54(2935), .W42TO55(13698), .W42TO56(3274), .W42TO57(-1641), .W42TO58(-10049), .W42TO59(19006), .W42TO60(221), .W42TO61(4064), .W42TO62(178), .W42TO63(-4249), .W42TO64(-9328), .W42TO65(1783), .W42TO66(-16119), .W42TO67(-7632), .W42TO68(21019), .W42TO69(-867), .W42TO70(1109), .W42TO71(-8213), .W42TO72(9651), .W42TO73(10524), .W42TO74(-10140), .W42TO75(15551), .W42TO76(11878), .W42TO77(-10012), .W42TO78(17925), .W42TO79(-17727), .W42TO80(21487), .W42TO81(-2636), .W42TO82(-12497), .W42TO83(-19715), .W42TO84(2742), .W42TO85(9498), .W42TO86(-21682), .W42TO87(3446), .W42TO88(-3526), .W42TO89(-232), .W42TO90(3841), .W42TO91(-10977), .W42TO92(20534), .W42TO93(3672), .W42TO94(-15988), .W42TO95(10650), .W42TO96(-1003), .W42TO97(20001), .W42TO98(-640), .W42TO99(3180), .W43TO0(-1866), .W43TO1(-10290), .W43TO2(-14040), .W43TO3(12699), .W43TO4(685), .W43TO5(-6894), .W43TO6(17835), .W43TO7(16152), .W43TO8(19258), .W43TO9(-5418), .W43TO10(6361), .W43TO11(7029), .W43TO12(-6687), .W43TO13(-7988), .W43TO14(-8789), .W43TO15(10144), .W43TO16(-10709), .W43TO17(11988), .W43TO18(-15980), .W43TO19(261), .W43TO20(-8445), .W43TO21(3568), .W43TO22(-8384), .W43TO23(-3614), .W43TO24(-269), .W43TO25(-5384), .W43TO26(-2561), .W43TO27(14404), .W43TO28(14504), .W43TO29(10021), .W43TO30(-11615), .W43TO31(20322), .W43TO32(5635), .W43TO33(-11968), .W43TO34(-11095), .W43TO35(13602), .W43TO36(8536), .W43TO37(6965), .W43TO38(15199), .W43TO39(3117), .W43TO40(7932), .W43TO41(18667), .W43TO42(-12078), .W43TO43(-12009), .W43TO44(5289), .W43TO45(-8970), .W43TO46(9408), .W43TO47(264), .W43TO48(-1464), .W43TO49(-30602), .W43TO50(2438), .W43TO51(-9806), .W43TO52(-15079), .W43TO53(-1252), .W43TO54(252), .W43TO55(3171), .W43TO56(8775), .W43TO57(-4176), .W43TO58(284), .W43TO59(3752), .W43TO60(17846), .W43TO61(725), .W43TO62(6693), .W43TO63(4901), .W43TO64(10674), .W43TO65(2347), .W43TO66(6207), .W43TO67(7505), .W43TO68(11345), .W43TO69(6232), .W43TO70(-8582), .W43TO71(-26383), .W43TO72(16341), .W43TO73(-12961), .W43TO74(-19060), .W43TO75(-9674), .W43TO76(-7955), .W43TO77(-13002), .W43TO78(19208), .W43TO79(-12817), .W43TO80(4394), .W43TO81(-14425), .W43TO82(2709), .W43TO83(-26638), .W43TO84(5106), .W43TO85(-2090), .W43TO86(-13989), .W43TO87(491), .W43TO88(-941), .W43TO89(-4870), .W43TO90(13577), .W43TO91(-18337), .W43TO92(74), .W43TO93(19515), .W43TO94(2090), .W43TO95(21076), .W43TO96(-715), .W43TO97(-10702), .W43TO98(9521), .W43TO99(7628), .W44TO0(-6605), .W44TO1(15506), .W44TO2(11111), .W44TO3(-17014), .W44TO4(-23158), .W44TO5(-7881), .W44TO6(-4397), .W44TO7(14527), .W44TO8(16655), .W44TO9(17171), .W44TO10(2063), .W44TO11(-387), .W44TO12(17316), .W44TO13(-6877), .W44TO14(11964), .W44TO15(3505), .W44TO16(-16573), .W44TO17(20809), .W44TO18(18739), .W44TO19(11537), .W44TO20(3965), .W44TO21(21066), .W44TO22(7461), .W44TO23(2472), .W44TO24(-3675), .W44TO25(-260), .W44TO26(8856), .W44TO27(-10237), .W44TO28(-12666), .W44TO29(-5707), .W44TO30(10765), .W44TO31(17030), .W44TO32(-12156), .W44TO33(-6227), .W44TO34(14919), .W44TO35(17076), .W44TO36(14084), .W44TO37(5944), .W44TO38(8172), .W44TO39(-5585), .W44TO40(6688), .W44TO41(-19227), .W44TO42(-17355), .W44TO43(-14727), .W44TO44(11974), .W44TO45(697), .W44TO46(-11697), .W44TO47(-3673), .W44TO48(-8749), .W44TO49(8612), .W44TO50(3361), .W44TO51(-6508), .W44TO52(-20274), .W44TO53(-5663), .W44TO54(-11627), .W44TO55(-503), .W44TO56(19059), .W44TO57(-16765), .W44TO58(5648), .W44TO59(-4041), .W44TO60(-4080), .W44TO61(13622), .W44TO62(-8356), .W44TO63(-2935), .W44TO64(-7192), .W44TO65(-5608), .W44TO66(-3826), .W44TO67(-5934), .W44TO68(1379), .W44TO69(-9818), .W44TO70(3325), .W44TO71(-3081), .W44TO72(15585), .W44TO73(7718), .W44TO74(-3216), .W44TO75(-1999), .W44TO76(6342), .W44TO77(655), .W44TO78(3223), .W44TO79(6232), .W44TO80(14618), .W44TO81(1652), .W44TO82(4742), .W44TO83(1041), .W44TO84(20437), .W44TO85(-6052), .W44TO86(12923), .W44TO87(2792), .W44TO88(-13711), .W44TO89(-13799), .W44TO90(-1842), .W44TO91(-10341), .W44TO92(-4438), .W44TO93(2989), .W44TO94(-14224), .W44TO95(22513), .W44TO96(7683), .W44TO97(-22233), .W44TO98(1336), .W44TO99(-8386), .W45TO0(-7360), .W45TO1(-7950), .W45TO2(-827), .W45TO3(10775), .W45TO4(-5439), .W45TO5(13352), .W45TO6(12330), .W45TO7(13514), .W45TO8(-3033), .W45TO9(-716), .W45TO10(8794), .W45TO11(-8184), .W45TO12(1424), .W45TO13(3866), .W45TO14(-15534), .W45TO15(14872), .W45TO16(1019), .W45TO17(-3513), .W45TO18(-13115), .W45TO19(-8989), .W45TO20(-9355), .W45TO21(1153), .W45TO22(10990), .W45TO23(-13812), .W45TO24(-1161), .W45TO25(22860), .W45TO26(8879), .W45TO27(-1180), .W45TO28(804), .W45TO29(15634), .W45TO30(20288), .W45TO31(14370), .W45TO32(22383), .W45TO33(18694), .W45TO34(9835), .W45TO35(-17361), .W45TO36(-12773), .W45TO37(-15198), .W45TO38(19978), .W45TO39(-3817), .W45TO40(5697), .W45TO41(17125), .W45TO42(-7554), .W45TO43(-8023), .W45TO44(13279), .W45TO45(4929), .W45TO46(-8651), .W45TO47(-8966), .W45TO48(-19874), .W45TO49(13865), .W45TO50(3781), .W45TO51(20906), .W45TO52(-683), .W45TO53(-3385), .W45TO54(-7870), .W45TO55(-9756), .W45TO56(-13152), .W45TO57(-19651), .W45TO58(-15206), .W45TO59(-5522), .W45TO60(-11572), .W45TO61(-285), .W45TO62(-3790), .W45TO63(5820), .W45TO64(-3876), .W45TO65(4850), .W45TO66(-5478), .W45TO67(-7666), .W45TO68(15088), .W45TO69(2916), .W45TO70(8517), .W45TO71(9606), .W45TO72(14706), .W45TO73(2120), .W45TO74(6014), .W45TO75(969), .W45TO76(8117), .W45TO77(2004), .W45TO78(-19184), .W45TO79(-3226), .W45TO80(8625), .W45TO81(-5296), .W45TO82(6951), .W45TO83(-11076), .W45TO84(-19906), .W45TO85(-1718), .W45TO86(7945), .W45TO87(20205), .W45TO88(-478), .W45TO89(-16619), .W45TO90(4328), .W45TO91(3511), .W45TO92(-11673), .W45TO93(18011), .W45TO94(9609), .W45TO95(-11459), .W45TO96(1066), .W45TO97(-7554), .W45TO98(-18590), .W45TO99(9748), .W46TO0(5977), .W46TO1(13019), .W46TO2(10689), .W46TO3(-5639), .W46TO4(-5773), .W46TO5(-2861), .W46TO6(6207), .W46TO7(-10393), .W46TO8(11246), .W46TO9(7351), .W46TO10(-15090), .W46TO11(6253), .W46TO12(-7798), .W46TO13(12859), .W46TO14(14843), .W46TO15(3380), .W46TO16(-12632), .W46TO17(-25254), .W46TO18(7258), .W46TO19(-13211), .W46TO20(6400), .W46TO21(-10423), .W46TO22(-7109), .W46TO23(19038), .W46TO24(14313), .W46TO25(-15092), .W46TO26(-12169), .W46TO27(8444), .W46TO28(-3843), .W46TO29(-7317), .W46TO30(15754), .W46TO31(-4137), .W46TO32(-10888), .W46TO33(17058), .W46TO34(5114), .W46TO35(18365), .W46TO36(-5277), .W46TO37(-14453), .W46TO38(-16676), .W46TO39(16745), .W46TO40(2300), .W46TO41(6155), .W46TO42(-16547), .W46TO43(10880), .W46TO44(10496), .W46TO45(2647), .W46TO46(-11250), .W46TO47(-8275), .W46TO48(-11014), .W46TO49(18224), .W46TO50(1497), .W46TO51(-1777), .W46TO52(-11596), .W46TO53(5959), .W46TO54(-2019), .W46TO55(15339), .W46TO56(9479), .W46TO57(-17710), .W46TO58(-6398), .W46TO59(-4728), .W46TO60(-7080), .W46TO61(-8980), .W46TO62(12686), .W46TO63(-4904), .W46TO64(10252), .W46TO65(-523), .W46TO66(12205), .W46TO67(4406), .W46TO68(5008), .W46TO69(-13074), .W46TO70(1429), .W46TO71(13233), .W46TO72(-2105), .W46TO73(-15731), .W46TO74(-3754), .W46TO75(-4177), .W46TO76(8069), .W46TO77(-19121), .W46TO78(3847), .W46TO79(19751), .W46TO80(-7261), .W46TO81(12936), .W46TO82(-9667), .W46TO83(-8525), .W46TO84(1326), .W46TO85(12117), .W46TO86(-20), .W46TO87(2075), .W46TO88(3600), .W46TO89(5817), .W46TO90(7552), .W46TO91(-9573), .W46TO92(11078), .W46TO93(6479), .W46TO94(258), .W46TO95(15048), .W46TO96(12895), .W46TO97(3864), .W46TO98(6670), .W46TO99(-13702), .W47TO0(-1991), .W47TO1(4490), .W47TO2(-17594), .W47TO3(15756), .W47TO4(-15065), .W47TO5(17011), .W47TO6(14645), .W47TO7(8908), .W47TO8(18089), .W47TO9(2726), .W47TO10(2848), .W47TO11(-15301), .W47TO12(-2308), .W47TO13(-16200), .W47TO14(6219), .W47TO15(-11764), .W47TO16(-17181), .W47TO17(3081), .W47TO18(3709), .W47TO19(17230), .W47TO20(-17141), .W47TO21(-9704), .W47TO22(17440), .W47TO23(16639), .W47TO24(-12042), .W47TO25(3166), .W47TO26(-6899), .W47TO27(-13785), .W47TO28(-3000), .W47TO29(-465), .W47TO30(5421), .W47TO31(10998), .W47TO32(5466), .W47TO33(9545), .W47TO34(7696), .W47TO35(4010), .W47TO36(8195), .W47TO37(9045), .W47TO38(-9862), .W47TO39(14566), .W47TO40(594), .W47TO41(-16013), .W47TO42(4853), .W47TO43(18014), .W47TO44(-1225), .W47TO45(19072), .W47TO46(-1828), .W47TO47(17409), .W47TO48(-18549), .W47TO49(-2422), .W47TO50(18437), .W47TO51(14797), .W47TO52(5238), .W47TO53(-7396), .W47TO54(15533), .W47TO55(-7571), .W47TO56(11160), .W47TO57(-5287), .W47TO58(5320), .W47TO59(1972), .W47TO60(-5566), .W47TO61(3804), .W47TO62(13202), .W47TO63(17559), .W47TO64(-13405), .W47TO65(6781), .W47TO66(-15900), .W47TO67(-4578), .W47TO68(-10047), .W47TO69(-16868), .W47TO70(-7825), .W47TO71(-4731), .W47TO72(7910), .W47TO73(8140), .W47TO74(13971), .W47TO75(1176), .W47TO76(18132), .W47TO77(16389), .W47TO78(-17561), .W47TO79(-932), .W47TO80(11415), .W47TO81(-6750), .W47TO82(-3196), .W47TO83(-15277), .W47TO84(-2329), .W47TO85(-6541), .W47TO86(4461), .W47TO87(-4612), .W47TO88(-5577), .W47TO89(2911), .W47TO90(-10530), .W47TO91(18884), .W47TO92(10593), .W47TO93(14432), .W47TO94(10233), .W47TO95(16304), .W47TO96(-17714), .W47TO97(7293), .W47TO98(-3156), .W47TO99(-17901), .W48TO0(3508), .W48TO1(18326), .W48TO2(-15881), .W48TO3(1797), .W48TO4(6703), .W48TO5(-18687), .W48TO6(18270), .W48TO7(1147), .W48TO8(-3538), .W48TO9(-5444), .W48TO10(9939), .W48TO11(-9136), .W48TO12(-12855), .W48TO13(10673), .W48TO14(-8303), .W48TO15(3105), .W48TO16(-6580), .W48TO17(13532), .W48TO18(5366), .W48TO19(-8847), .W48TO20(-17371), .W48TO21(-9841), .W48TO22(10708), .W48TO23(-6326), .W48TO24(14954), .W48TO25(-18613), .W48TO26(-8009), .W48TO27(-12894), .W48TO28(-9101), .W48TO29(-3294), .W48TO30(3805), .W48TO31(-9702), .W48TO32(-12391), .W48TO33(-6638), .W48TO34(538), .W48TO35(-12308), .W48TO36(5378), .W48TO37(-18676), .W48TO38(15765), .W48TO39(7959), .W48TO40(-16890), .W48TO41(18530), .W48TO42(18951), .W48TO43(-6988), .W48TO44(-14861), .W48TO45(-15249), .W48TO46(16954), .W48TO47(8304), .W48TO48(2463), .W48TO49(-13998), .W48TO50(-10560), .W48TO51(-13906), .W48TO52(-13600), .W48TO53(17183), .W48TO54(18236), .W48TO55(11720), .W48TO56(938), .W48TO57(12205), .W48TO58(-11850), .W48TO59(-2622), .W48TO60(-1098), .W48TO61(18067), .W48TO62(16861), .W48TO63(-15301), .W48TO64(-6565), .W48TO65(-5967), .W48TO66(-13646), .W48TO67(18250), .W48TO68(14211), .W48TO69(-2805), .W48TO70(7140), .W48TO71(1245), .W48TO72(-8815), .W48TO73(-9891), .W48TO74(-2329), .W48TO75(-2345), .W48TO76(3524), .W48TO77(-6537), .W48TO78(8901), .W48TO79(10763), .W48TO80(17543), .W48TO81(-10337), .W48TO82(2655), .W48TO83(-2882), .W48TO84(-13577), .W48TO85(12653), .W48TO86(-15883), .W48TO87(-9872), .W48TO88(4209), .W48TO89(3429), .W48TO90(15764), .W48TO91(15374), .W48TO92(11765), .W48TO93(-860), .W48TO94(10299), .W48TO95(17577), .W48TO96(16575), .W48TO97(-5691), .W48TO98(-4616), .W48TO99(-19099), .W49TO0(13445), .W49TO1(11239), .W49TO2(404), .W49TO3(-18433), .W49TO4(-18415), .W49TO5(12154), .W49TO6(-13926), .W49TO7(987), .W49TO8(11412), .W49TO9(1329), .W49TO10(-3413), .W49TO11(-18277), .W49TO12(3782), .W49TO13(12256), .W49TO14(14771), .W49TO15(13729), .W49TO16(-10702), .W49TO17(-14097), .W49TO18(-10466), .W49TO19(-9898), .W49TO20(6870), .W49TO21(8917), .W49TO22(16056), .W49TO23(-6383), .W49TO24(-9496), .W49TO25(18365), .W49TO26(11025), .W49TO27(-18828), .W49TO28(-6762), .W49TO29(-11666), .W49TO30(14673), .W49TO31(2887), .W49TO32(11199), .W49TO33(-1727), .W49TO34(-754), .W49TO35(16964), .W49TO36(7482), .W49TO37(-610), .W49TO38(-16223), .W49TO39(-8373), .W49TO40(-13738), .W49TO41(12951), .W49TO42(18589), .W49TO43(8733), .W49TO44(18604), .W49TO45(-5523), .W49TO46(-12157), .W49TO47(5524), .W49TO48(-7404), .W49TO49(-5686), .W49TO50(6685), .W49TO51(4185), .W49TO52(2907), .W49TO53(-18521), .W49TO54(-6629), .W49TO55(7566), .W49TO56(-13035), .W49TO57(-13719), .W49TO58(14022), .W49TO59(-13336), .W49TO60(-6603), .W49TO61(-8620), .W49TO62(-17027), .W49TO63(10618), .W49TO64(15705), .W49TO65(-7603), .W49TO66(1724), .W49TO67(-3116), .W49TO68(-13649), .W49TO69(14101), .W49TO70(12917), .W49TO71(16148), .W49TO72(-371), .W49TO73(-8489), .W49TO74(11998), .W49TO75(11901), .W49TO76(18027), .W49TO77(15535), .W49TO78(-118), .W49TO79(16863), .W49TO80(17412), .W49TO81(-7133), .W49TO82(-15724), .W49TO83(-15250), .W49TO84(11512), .W49TO85(6796), .W49TO86(-11701), .W49TO87(-11570), .W49TO88(10170), .W49TO89(-14022), .W49TO90(-9668), .W49TO91(6888), .W49TO92(-10637), .W49TO93(-8916), .W49TO94(-11698), .W49TO95(10154), .W49TO96(11475), .W49TO97(12405), .W49TO98(-9007), .W49TO99(-4862), .W50TO0(-572), .W50TO1(10807), .W50TO2(-1623), .W50TO3(-2645), .W50TO4(-7687), .W50TO5(-2573), .W50TO6(-3636), .W50TO7(2937), .W50TO8(-13754), .W50TO9(1479), .W50TO10(10055), .W50TO11(-17325), .W50TO12(-5209), .W50TO13(3121), .W50TO14(14968), .W50TO15(-8132), .W50TO16(-901), .W50TO17(-2231), .W50TO18(-18241), .W50TO19(1343), .W50TO20(2744), .W50TO21(-14712), .W50TO22(-16650), .W50TO23(-13512), .W50TO24(2993), .W50TO25(-3850), .W50TO26(-13960), .W50TO27(2016), .W50TO28(-16093), .W50TO29(760), .W50TO30(13552), .W50TO31(3322), .W50TO32(-14834), .W50TO33(-13084), .W50TO34(685), .W50TO35(6638), .W50TO36(13584), .W50TO37(20600), .W50TO38(20735), .W50TO39(-20963), .W50TO40(10847), .W50TO41(529), .W50TO42(-1010), .W50TO43(-5798), .W50TO44(-5409), .W50TO45(1457), .W50TO46(7578), .W50TO47(627), .W50TO48(-13404), .W50TO49(-10191), .W50TO50(-2880), .W50TO51(19467), .W50TO52(-13988), .W50TO53(-16487), .W50TO54(6576), .W50TO55(-16688), .W50TO56(9506), .W50TO57(15192), .W50TO58(-4813), .W50TO59(179), .W50TO60(-15103), .W50TO61(19772), .W50TO62(-7511), .W50TO63(7969), .W50TO64(-778), .W50TO65(-18995), .W50TO66(3437), .W50TO67(10106), .W50TO68(-11702), .W50TO69(6034), .W50TO70(17420), .W50TO71(-20977), .W50TO72(-5681), .W50TO73(-3516), .W50TO74(-17716), .W50TO75(-4993), .W50TO76(-108), .W50TO77(19357), .W50TO78(-10374), .W50TO79(-13729), .W50TO80(20308), .W50TO81(11892), .W50TO82(2754), .W50TO83(-2010), .W50TO84(-9744), .W50TO85(-16004), .W50TO86(-2391), .W50TO87(18184), .W50TO88(9895), .W50TO89(-7234), .W50TO90(-13806), .W50TO91(769), .W50TO92(-2032), .W50TO93(6541), .W50TO94(-21494), .W50TO95(12076), .W50TO96(-9368), .W50TO97(439), .W50TO98(12520), .W50TO99(11584), .W51TO0(-2522), .W51TO1(11653), .W51TO2(13875), .W51TO3(6328), .W51TO4(17377), .W51TO5(1460), .W51TO6(-199), .W51TO7(-4500), .W51TO8(11285), .W51TO9(4275), .W51TO10(4973), .W51TO11(16645), .W51TO12(-8993), .W51TO13(-4659), .W51TO14(886), .W51TO15(8225), .W51TO16(894), .W51TO17(10229), .W51TO18(15080), .W51TO19(8368), .W51TO20(3606), .W51TO21(-857), .W51TO22(-9069), .W51TO23(-10870), .W51TO24(2190), .W51TO25(-16107), .W51TO26(-732), .W51TO27(-15536), .W51TO28(3433), .W51TO29(-18617), .W51TO30(13591), .W51TO31(-2247), .W51TO32(11787), .W51TO33(-747), .W51TO34(8679), .W51TO35(16779), .W51TO36(10539), .W51TO37(15070), .W51TO38(9075), .W51TO39(-9878), .W51TO40(-17327), .W51TO41(-11157), .W51TO42(2241), .W51TO43(-2830), .W51TO44(4327), .W51TO45(9877), .W51TO46(12808), .W51TO47(-15890), .W51TO48(-13562), .W51TO49(-25994), .W51TO50(-6405), .W51TO51(-1923), .W51TO52(12444), .W51TO53(20), .W51TO54(-9221), .W51TO55(5264), .W51TO56(2534), .W51TO57(-14726), .W51TO58(16818), .W51TO59(17347), .W51TO60(1130), .W51TO61(-14673), .W51TO62(-19337), .W51TO63(14717), .W51TO64(17301), .W51TO65(-15225), .W51TO66(-15575), .W51TO67(3420), .W51TO68(19906), .W51TO69(-10181), .W51TO70(82), .W51TO71(1311), .W51TO72(10213), .W51TO73(-10454), .W51TO74(-10722), .W51TO75(9012), .W51TO76(-15490), .W51TO77(-3930), .W51TO78(3997), .W51TO79(-15751), .W51TO80(1230), .W51TO81(834), .W51TO82(-2740), .W51TO83(7829), .W51TO84(-15107), .W51TO85(-2090), .W51TO86(5475), .W51TO87(-8498), .W51TO88(11083), .W51TO89(16029), .W51TO90(18946), .W51TO91(-8924), .W51TO92(10671), .W51TO93(12905), .W51TO94(-8712), .W51TO95(8422), .W51TO96(14529), .W51TO97(-3291), .W51TO98(-2353), .W51TO99(14501), .W52TO0(-653), .W52TO1(19241), .W52TO2(13141), .W52TO3(474), .W52TO4(1170), .W52TO5(-5120), .W52TO6(-1200), .W52TO7(-13941), .W52TO8(-11168), .W52TO9(-5276), .W52TO10(7237), .W52TO11(2705), .W52TO12(1129), .W52TO13(-328), .W52TO14(14002), .W52TO15(5262), .W52TO16(-4155), .W52TO17(-717), .W52TO18(17452), .W52TO19(-10110), .W52TO20(-1346), .W52TO21(-8005), .W52TO22(-12150), .W52TO23(-5504), .W52TO24(7575), .W52TO25(-13463), .W52TO26(23), .W52TO27(5854), .W52TO28(-1332), .W52TO29(9523), .W52TO30(-7397), .W52TO31(8122), .W52TO32(-7077), .W52TO33(-8332), .W52TO34(-9091), .W52TO35(1031), .W52TO36(14290), .W52TO37(-3557), .W52TO38(19811), .W52TO39(-874), .W52TO40(4792), .W52TO41(934), .W52TO42(8601), .W52TO43(23490), .W52TO44(6790), .W52TO45(6433), .W52TO46(-8820), .W52TO47(-22750), .W52TO48(12450), .W52TO49(4641), .W52TO50(-4618), .W52TO51(-673), .W52TO52(-3376), .W52TO53(6257), .W52TO54(-15763), .W52TO55(-10723), .W52TO56(-1234), .W52TO57(11041), .W52TO58(11733), .W52TO59(-1219), .W52TO60(971), .W52TO61(-9145), .W52TO62(4616), .W52TO63(-5574), .W52TO64(5411), .W52TO65(14854), .W52TO66(-1950), .W52TO67(24974), .W52TO68(-13190), .W52TO69(2410), .W52TO70(-13256), .W52TO71(4934), .W52TO72(-8062), .W52TO73(5687), .W52TO74(9774), .W52TO75(10157), .W52TO76(20535), .W52TO77(-2062), .W52TO78(14826), .W52TO79(-11254), .W52TO80(-485), .W52TO81(-1679), .W52TO82(6574), .W52TO83(11323), .W52TO84(-5799), .W52TO85(-1087), .W52TO86(-6741), .W52TO87(-6479), .W52TO88(-15385), .W52TO89(6366), .W52TO90(2640), .W52TO91(-8042), .W52TO92(19424), .W52TO93(-4255), .W52TO94(4507), .W52TO95(14268), .W52TO96(-1072), .W52TO97(-8147), .W52TO98(-537), .W52TO99(9356), .W53TO0(-16840), .W53TO1(7514), .W53TO2(-2529), .W53TO3(-14000), .W53TO4(21790), .W53TO5(-15483), .W53TO6(12611), .W53TO7(-22727), .W53TO8(-12541), .W53TO9(-489), .W53TO10(4301), .W53TO11(-4209), .W53TO12(3685), .W53TO13(12932), .W53TO14(-8302), .W53TO15(981), .W53TO16(-16780), .W53TO17(-9136), .W53TO18(-4197), .W53TO19(26043), .W53TO20(7307), .W53TO21(5844), .W53TO22(5535), .W53TO23(15318), .W53TO24(-7555), .W53TO25(-11063), .W53TO26(-13312), .W53TO27(1050), .W53TO28(-8853), .W53TO29(-18344), .W53TO30(-8459), .W53TO31(-16084), .W53TO32(16781), .W53TO33(-6142), .W53TO34(-4410), .W53TO35(16958), .W53TO36(-13619), .W53TO37(7194), .W53TO38(-13677), .W53TO39(-17179), .W53TO40(-5416), .W53TO41(21250), .W53TO42(6165), .W53TO43(-9399), .W53TO44(-6694), .W53TO45(-10701), .W53TO46(-1392), .W53TO47(6966), .W53TO48(9797), .W53TO49(7189), .W53TO50(-13940), .W53TO51(13976), .W53TO52(-7012), .W53TO53(17505), .W53TO54(19159), .W53TO55(-6865), .W53TO56(9107), .W53TO57(-11981), .W53TO58(3529), .W53TO59(16665), .W53TO60(-1454), .W53TO61(155), .W53TO62(-6776), .W53TO63(-9422), .W53TO64(12584), .W53TO65(-6136), .W53TO66(-19767), .W53TO67(18043), .W53TO68(-5022), .W53TO69(16459), .W53TO70(6414), .W53TO71(13257), .W53TO72(9109), .W53TO73(-11065), .W53TO74(-185), .W53TO75(-7394), .W53TO76(15487), .W53TO77(-11507), .W53TO78(10910), .W53TO79(-2371), .W53TO80(422), .W53TO81(-12625), .W53TO82(19324), .W53TO83(1552), .W53TO84(433), .W53TO85(-12680), .W53TO86(-8192), .W53TO87(-3125), .W53TO88(8204), .W53TO89(20928), .W53TO90(12794), .W53TO91(2758), .W53TO92(10047), .W53TO93(-3540), .W53TO94(-12757), .W53TO95(13537), .W53TO96(-3633), .W53TO97(-13711), .W53TO98(20359), .W53TO99(-18106), .W54TO0(12417), .W54TO1(-5499), .W54TO2(14102), .W54TO3(13522), .W54TO4(15379), .W54TO5(6874), .W54TO6(-16173), .W54TO7(11569), .W54TO8(-17801), .W54TO9(-7684), .W54TO10(-15525), .W54TO11(7972), .W54TO12(-15639), .W54TO13(-5735), .W54TO14(-15198), .W54TO15(-3176), .W54TO16(9980), .W54TO17(3267), .W54TO18(14449), .W54TO19(14945), .W54TO20(-7004), .W54TO21(-4401), .W54TO22(6378), .W54TO23(12186), .W54TO24(-444), .W54TO25(1984), .W54TO26(9214), .W54TO27(16590), .W54TO28(-947), .W54TO29(12182), .W54TO30(-9468), .W54TO31(12109), .W54TO32(-10478), .W54TO33(-4419), .W54TO34(15277), .W54TO35(14580), .W54TO36(5325), .W54TO37(-4883), .W54TO38(-3399), .W54TO39(-12656), .W54TO40(6962), .W54TO41(-6945), .W54TO42(8864), .W54TO43(5976), .W54TO44(9880), .W54TO45(-10651), .W54TO46(3789), .W54TO47(-9113), .W54TO48(13621), .W54TO49(-11104), .W54TO50(1338), .W54TO51(5250), .W54TO52(8178), .W54TO53(10697), .W54TO54(-1772), .W54TO55(113), .W54TO56(16576), .W54TO57(7836), .W54TO58(909), .W54TO59(14164), .W54TO60(904), .W54TO61(-6375), .W54TO62(-17744), .W54TO63(15776), .W54TO64(6906), .W54TO65(-13788), .W54TO66(6623), .W54TO67(8429), .W54TO68(12637), .W54TO69(7993), .W54TO70(11889), .W54TO71(13139), .W54TO72(15931), .W54TO73(1133), .W54TO74(-10571), .W54TO75(12922), .W54TO76(2779), .W54TO77(6844), .W54TO78(-11790), .W54TO79(-7498), .W54TO80(-8967), .W54TO81(5137), .W54TO82(2711), .W54TO83(6148), .W54TO84(-15733), .W54TO85(3581), .W54TO86(17859), .W54TO87(10453), .W54TO88(-1399), .W54TO89(21119), .W54TO90(-3872), .W54TO91(-1476), .W54TO92(-6432), .W54TO93(-13914), .W54TO94(5045), .W54TO95(-13520), .W54TO96(-7659), .W54TO97(2036), .W54TO98(-12693), .W54TO99(12511), .W55TO0(9300), .W55TO1(-4627), .W55TO2(16774), .W55TO3(-12397), .W55TO4(11309), .W55TO5(-14447), .W55TO6(-18178), .W55TO7(-7907), .W55TO8(2542), .W55TO9(-430), .W55TO10(-14738), .W55TO11(-6239), .W55TO12(4205), .W55TO13(-3210), .W55TO14(-17764), .W55TO15(-18067), .W55TO16(-17515), .W55TO17(13245), .W55TO18(17173), .W55TO19(17609), .W55TO20(4935), .W55TO21(-6879), .W55TO22(14630), .W55TO23(2350), .W55TO24(-2731), .W55TO25(1563), .W55TO26(10043), .W55TO27(-11456), .W55TO28(-3606), .W55TO29(15740), .W55TO30(-16663), .W55TO31(16438), .W55TO32(-5329), .W55TO33(-17356), .W55TO34(-9852), .W55TO35(-5408), .W55TO36(9868), .W55TO37(-9872), .W55TO38(-5679), .W55TO39(11503), .W55TO40(-2069), .W55TO41(4043), .W55TO42(17675), .W55TO43(-7606), .W55TO44(16254), .W55TO45(2956), .W55TO46(-3465), .W55TO47(-1563), .W55TO48(3721), .W55TO49(-18809), .W55TO50(3802), .W55TO51(12618), .W55TO52(-8429), .W55TO53(15977), .W55TO54(16347), .W55TO55(9287), .W55TO56(3768), .W55TO57(-7961), .W55TO58(6051), .W55TO59(17313), .W55TO60(11526), .W55TO61(12173), .W55TO62(-11422), .W55TO63(-4582), .W55TO64(9202), .W55TO65(715), .W55TO66(-13618), .W55TO67(-1366), .W55TO68(4036), .W55TO69(-8306), .W55TO70(17806), .W55TO71(5065), .W55TO72(18982), .W55TO73(8344), .W55TO74(-11655), .W55TO75(-10168), .W55TO76(-3387), .W55TO77(12583), .W55TO78(5285), .W55TO79(9909), .W55TO80(-6195), .W55TO81(14299), .W55TO82(-9176), .W55TO83(279), .W55TO84(4392), .W55TO85(-453), .W55TO86(10808), .W55TO87(-3211), .W55TO88(15628), .W55TO89(-2524), .W55TO90(-12237), .W55TO91(-15092), .W55TO92(4151), .W55TO93(-15887), .W55TO94(16085), .W55TO95(5335), .W55TO96(11926), .W55TO97(-13140), .W55TO98(-5252), .W55TO99(-1354), .W56TO0(1687), .W56TO1(6488), .W56TO2(-11988), .W56TO3(-8748), .W56TO4(13544), .W56TO5(3155), .W56TO6(-1147), .W56TO7(335), .W56TO8(-18684), .W56TO9(-10178), .W56TO10(4244), .W56TO11(-1053), .W56TO12(-7814), .W56TO13(10884), .W56TO14(-12100), .W56TO15(-2241), .W56TO16(1940), .W56TO17(-10095), .W56TO18(-8942), .W56TO19(18557), .W56TO20(-3754), .W56TO21(-11863), .W56TO22(-16504), .W56TO23(-17404), .W56TO24(14738), .W56TO25(-2015), .W56TO26(-9042), .W56TO27(3819), .W56TO28(-13809), .W56TO29(-119), .W56TO30(4542), .W56TO31(-319), .W56TO32(-9931), .W56TO33(-6459), .W56TO34(-5658), .W56TO35(6623), .W56TO36(-18944), .W56TO37(3193), .W56TO38(16081), .W56TO39(6317), .W56TO40(11073), .W56TO41(-12472), .W56TO42(-7617), .W56TO43(-2139), .W56TO44(16537), .W56TO45(-11097), .W56TO46(-5303), .W56TO47(5733), .W56TO48(13385), .W56TO49(-4318), .W56TO50(2674), .W56TO51(11897), .W56TO52(12772), .W56TO53(-12302), .W56TO54(17198), .W56TO55(-12483), .W56TO56(-13557), .W56TO57(10476), .W56TO58(-6092), .W56TO59(-4674), .W56TO60(7901), .W56TO61(11607), .W56TO62(-2832), .W56TO63(-16161), .W56TO64(3847), .W56TO65(15858), .W56TO66(7084), .W56TO67(-14178), .W56TO68(9801), .W56TO69(-16064), .W56TO70(-18822), .W56TO71(-12067), .W56TO72(-11443), .W56TO73(-14917), .W56TO74(13410), .W56TO75(-4365), .W56TO76(-13262), .W56TO77(-3038), .W56TO78(-3421), .W56TO79(7364), .W56TO80(-7240), .W56TO81(-1525), .W56TO82(-8561), .W56TO83(13724), .W56TO84(-10571), .W56TO85(2583), .W56TO86(1381), .W56TO87(18552), .W56TO88(10038), .W56TO89(-13086), .W56TO90(7775), .W56TO91(-5656), .W56TO92(154), .W56TO93(-2722), .W56TO94(-17637), .W56TO95(887), .W56TO96(-5288), .W56TO97(-3296), .W56TO98(17270), .W56TO99(138), .W57TO0(-7582), .W57TO1(744), .W57TO2(9355), .W57TO3(-3938), .W57TO4(-11796), .W57TO5(2336), .W57TO6(-12979), .W57TO7(17678), .W57TO8(-12894), .W57TO9(17262), .W57TO10(5924), .W57TO11(-6129), .W57TO12(-889), .W57TO13(-9750), .W57TO14(-16515), .W57TO15(-12448), .W57TO16(-12291), .W57TO17(-15475), .W57TO18(-14417), .W57TO19(-1781), .W57TO20(12682), .W57TO21(-7245), .W57TO22(-6553), .W57TO23(16385), .W57TO24(-6942), .W57TO25(10559), .W57TO26(-5888), .W57TO27(-5327), .W57TO28(-18082), .W57TO29(8357), .W57TO30(-10070), .W57TO31(12925), .W57TO32(-2773), .W57TO33(9428), .W57TO34(-13290), .W57TO35(-9893), .W57TO36(-10154), .W57TO37(7886), .W57TO38(3416), .W57TO39(-15127), .W57TO40(10209), .W57TO41(-9290), .W57TO42(1668), .W57TO43(3544), .W57TO44(-9244), .W57TO45(-2197), .W57TO46(15671), .W57TO47(3922), .W57TO48(-8222), .W57TO49(7405), .W57TO50(-73), .W57TO51(14655), .W57TO52(3329), .W57TO53(-15636), .W57TO54(4045), .W57TO55(-1368), .W57TO56(-1138), .W57TO57(-9304), .W57TO58(-11159), .W57TO59(15243), .W57TO60(-16305), .W57TO61(6492), .W57TO62(12099), .W57TO63(-10081), .W57TO64(15037), .W57TO65(12979), .W57TO66(-6630), .W57TO67(11676), .W57TO68(3549), .W57TO69(18814), .W57TO70(18180), .W57TO71(-6994), .W57TO72(3706), .W57TO73(-15488), .W57TO74(-18262), .W57TO75(-11883), .W57TO76(18719), .W57TO77(4415), .W57TO78(12262), .W57TO79(-4661), .W57TO80(1268), .W57TO81(7706), .W57TO82(12779), .W57TO83(11081), .W57TO84(-8660), .W57TO85(9940), .W57TO86(-4881), .W57TO87(-12151), .W57TO88(-2214), .W57TO89(-14376), .W57TO90(-15123), .W57TO91(14392), .W57TO92(-11365), .W57TO93(-16473), .W57TO94(-6250), .W57TO95(-16346), .W57TO96(-7338), .W57TO97(-5650), .W57TO98(-6822), .W57TO99(12862), .W58TO0(-3108), .W58TO1(-13338), .W58TO2(-13505), .W58TO3(2662), .W58TO4(12450), .W58TO5(20784), .W58TO6(-15678), .W58TO7(-5978), .W58TO8(2103), .W58TO9(18687), .W58TO10(18977), .W58TO11(13490), .W58TO12(-3975), .W58TO13(-3970), .W58TO14(17465), .W58TO15(-814), .W58TO16(3080), .W58TO17(-7617), .W58TO18(3766), .W58TO19(13941), .W58TO20(11787), .W58TO21(-15243), .W58TO22(6984), .W58TO23(-19682), .W58TO24(22471), .W58TO25(4939), .W58TO26(-2194), .W58TO27(-3247), .W58TO28(-3050), .W58TO29(-4303), .W58TO30(-14092), .W58TO31(-20786), .W58TO32(11735), .W58TO33(2828), .W58TO34(2128), .W58TO35(-877), .W58TO36(2153), .W58TO37(-12027), .W58TO38(-12829), .W58TO39(11284), .W58TO40(-19059), .W58TO41(-3845), .W58TO42(-15519), .W58TO43(-4835), .W58TO44(-9888), .W58TO45(-3571), .W58TO46(9263), .W58TO47(2473), .W58TO48(-16789), .W58TO49(-1650), .W58TO50(11784), .W58TO51(17695), .W58TO52(-5827), .W58TO53(4155), .W58TO54(-7827), .W58TO55(-5828), .W58TO56(15221), .W58TO57(-14906), .W58TO58(-12379), .W58TO59(4578), .W58TO60(4831), .W58TO61(-8673), .W58TO62(-17295), .W58TO63(3271), .W58TO64(-9028), .W58TO65(-10094), .W58TO66(-5715), .W58TO67(946), .W58TO68(2955), .W58TO69(-15249), .W58TO70(-12207), .W58TO71(-19761), .W58TO72(-9585), .W58TO73(13090), .W58TO74(-17236), .W58TO75(11443), .W58TO76(8431), .W58TO77(12374), .W58TO78(3996), .W58TO79(18519), .W58TO80(-14504), .W58TO81(18148), .W58TO82(9752), .W58TO83(17206), .W58TO84(-10102), .W58TO85(-17414), .W58TO86(-15073), .W58TO87(-926), .W58TO88(-9745), .W58TO89(21450), .W58TO90(-1106), .W58TO91(2981), .W58TO92(-11986), .W58TO93(1235), .W58TO94(5785), .W58TO95(-1143), .W58TO96(-15214), .W58TO97(11295), .W58TO98(-11916), .W58TO99(17014), .W59TO0(14814), .W59TO1(-16862), .W59TO2(-3478), .W59TO3(-10415), .W59TO4(-8393), .W59TO5(4340), .W59TO6(14980), .W59TO7(-20428), .W59TO8(-1687), .W59TO9(1653), .W59TO10(2585), .W59TO11(1613), .W59TO12(17406), .W59TO13(12603), .W59TO14(15985), .W59TO15(-4643), .W59TO16(-8109), .W59TO17(804), .W59TO18(-3721), .W59TO19(903), .W59TO20(11346), .W59TO21(6176), .W59TO22(8668), .W59TO23(3688), .W59TO24(15293), .W59TO25(-14648), .W59TO26(-11176), .W59TO27(-9291), .W59TO28(13238), .W59TO29(5017), .W59TO30(-13316), .W59TO31(14760), .W59TO32(731), .W59TO33(-2181), .W59TO34(-20040), .W59TO35(7299), .W59TO36(-9221), .W59TO37(20538), .W59TO38(-2969), .W59TO39(-20806), .W59TO40(-14936), .W59TO41(-3598), .W59TO42(-17250), .W59TO43(15582), .W59TO44(9218), .W59TO45(-19684), .W59TO46(-12583), .W59TO47(9542), .W59TO48(-12131), .W59TO49(14511), .W59TO50(918), .W59TO51(7036), .W59TO52(2664), .W59TO53(-2939), .W59TO54(-17068), .W59TO55(-17458), .W59TO56(6794), .W59TO57(14423), .W59TO58(-8708), .W59TO59(-9395), .W59TO60(-14208), .W59TO61(-3218), .W59TO62(7314), .W59TO63(7446), .W59TO64(-4460), .W59TO65(-17736), .W59TO66(-6586), .W59TO67(3874), .W59TO68(14), .W59TO69(8034), .W59TO70(9371), .W59TO71(6520), .W59TO72(2678), .W59TO73(10117), .W59TO74(11007), .W59TO75(-16519), .W59TO76(-4787), .W59TO77(-6242), .W59TO78(1416), .W59TO79(-13028), .W59TO80(-8513), .W59TO81(-2911), .W59TO82(3627), .W59TO83(175), .W59TO84(1459), .W59TO85(4250), .W59TO86(-9353), .W59TO87(1722), .W59TO88(-4117), .W59TO89(22623), .W59TO90(5109), .W59TO91(-3176), .W59TO92(-1039), .W59TO93(8086), .W59TO94(10084), .W59TO95(-19157), .W59TO96(-18670), .W59TO97(2921), .W59TO98(-8714), .W59TO99(-1340), .W60TO0(-17600), .W60TO1(3378), .W60TO2(-8848), .W60TO3(-23071), .W60TO4(-480), .W60TO5(-3647), .W60TO6(6936), .W60TO7(-17204), .W60TO8(5544), .W60TO9(-2387), .W60TO10(18104), .W60TO11(17677), .W60TO12(-11781), .W60TO13(-5076), .W60TO14(-15758), .W60TO15(-16551), .W60TO16(2484), .W60TO17(-13495), .W60TO18(14749), .W60TO19(20127), .W60TO20(7588), .W60TO21(-3122), .W60TO22(-19614), .W60TO23(6217), .W60TO24(-7842), .W60TO25(-11097), .W60TO26(-21149), .W60TO27(-12575), .W60TO28(-14222), .W60TO29(-13642), .W60TO30(-9769), .W60TO31(-15072), .W60TO32(11806), .W60TO33(6817), .W60TO34(-2562), .W60TO35(-4121), .W60TO36(1978), .W60TO37(-12057), .W60TO38(7655), .W60TO39(4916), .W60TO40(5144), .W60TO41(5186), .W60TO42(-23721), .W60TO43(25059), .W60TO44(18310), .W60TO45(2006), .W60TO46(-4714), .W60TO47(-5432), .W60TO48(-13477), .W60TO49(4517), .W60TO50(-10512), .W60TO51(-7366), .W60TO52(18180), .W60TO53(14259), .W60TO54(252), .W60TO55(-4784), .W60TO56(16276), .W60TO57(-10893), .W60TO58(-16486), .W60TO59(-3397), .W60TO60(-4026), .W60TO61(-7274), .W60TO62(-8595), .W60TO63(-4410), .W60TO64(-8217), .W60TO65(-6268), .W60TO66(-19954), .W60TO67(13725), .W60TO68(-2998), .W60TO69(-1425), .W60TO70(9835), .W60TO71(-10664), .W60TO72(20835), .W60TO73(-13166), .W60TO74(-11647), .W60TO75(-18652), .W60TO76(-9054), .W60TO77(490), .W60TO78(-16637), .W60TO79(-5265), .W60TO80(4607), .W60TO81(5128), .W60TO82(5433), .W60TO83(-729), .W60TO84(-14394), .W60TO85(5203), .W60TO86(20838), .W60TO87(-9640), .W60TO88(13525), .W60TO89(-2975), .W60TO90(6794), .W60TO91(16662), .W60TO92(19686), .W60TO93(12352), .W60TO94(-22010), .W60TO95(2010), .W60TO96(7793), .W60TO97(-6386), .W60TO98(20405), .W60TO99(8591), .W61TO0(-14295), .W61TO1(15786), .W61TO2(2734), .W61TO3(-19487), .W61TO4(-7086), .W61TO5(-3103), .W61TO6(-5817), .W61TO7(-13289), .W61TO8(-6845), .W61TO9(8286), .W61TO10(-5537), .W61TO11(-14297), .W61TO12(-17398), .W61TO13(-1598), .W61TO14(-9425), .W61TO15(18674), .W61TO16(9705), .W61TO17(-11086), .W61TO18(180), .W61TO19(3589), .W61TO20(-8946), .W61TO21(-6991), .W61TO22(9530), .W61TO23(12912), .W61TO24(1133), .W61TO25(24167), .W61TO26(15804), .W61TO27(-18776), .W61TO28(-8059), .W61TO29(-15141), .W61TO30(18771), .W61TO31(4725), .W61TO32(20064), .W61TO33(-8658), .W61TO34(-2528), .W61TO35(-15144), .W61TO36(3229), .W61TO37(12542), .W61TO38(-5414), .W61TO39(-20795), .W61TO40(-11499), .W61TO41(642), .W61TO42(-14911), .W61TO43(12349), .W61TO44(10714), .W61TO45(-8373), .W61TO46(-274), .W61TO47(3095), .W61TO48(-2559), .W61TO49(499), .W61TO50(-6984), .W61TO51(-102), .W61TO52(19870), .W61TO53(-3937), .W61TO54(2602), .W61TO55(-219), .W61TO56(14501), .W61TO57(15303), .W61TO58(19594), .W61TO59(-10284), .W61TO60(-4554), .W61TO61(9700), .W61TO62(5636), .W61TO63(6454), .W61TO64(-12734), .W61TO65(-3104), .W61TO66(-11640), .W61TO67(17913), .W61TO68(-856), .W61TO69(4190), .W61TO70(3534), .W61TO71(-9979), .W61TO72(19967), .W61TO73(3444), .W61TO74(17035), .W61TO75(-9235), .W61TO76(12253), .W61TO77(-10553), .W61TO78(17015), .W61TO79(-434), .W61TO80(8601), .W61TO81(-8017), .W61TO82(23850), .W61TO83(9345), .W61TO84(13832), .W61TO85(14049), .W61TO86(-9081), .W61TO87(-21153), .W61TO88(-1632), .W61TO89(11202), .W61TO90(-2377), .W61TO91(11576), .W61TO92(-7081), .W61TO93(-3084), .W61TO94(8700), .W61TO95(9994), .W61TO96(-78), .W61TO97(-10389), .W61TO98(15978), .W61TO99(10540), .W62TO0(-5963), .W62TO1(-1033), .W62TO2(-13096), .W62TO3(16739), .W62TO4(15612), .W62TO5(-21492), .W62TO6(3989), .W62TO7(11689), .W62TO8(-15649), .W62TO9(-4547), .W62TO10(-8044), .W62TO11(-6434), .W62TO12(11530), .W62TO13(19562), .W62TO14(287), .W62TO15(13674), .W62TO16(-9489), .W62TO17(11182), .W62TO18(18788), .W62TO19(10643), .W62TO20(-17970), .W62TO21(-14559), .W62TO22(-16360), .W62TO23(11376), .W62TO24(8043), .W62TO25(19774), .W62TO26(3387), .W62TO27(-23), .W62TO28(-15285), .W62TO29(-5166), .W62TO30(-19340), .W62TO31(12948), .W62TO32(16849), .W62TO33(-5126), .W62TO34(9601), .W62TO35(3797), .W62TO36(-3853), .W62TO37(16057), .W62TO38(14885), .W62TO39(16323), .W62TO40(-12618), .W62TO41(168), .W62TO42(2867), .W62TO43(-7505), .W62TO44(6009), .W62TO45(-7010), .W62TO46(-16327), .W62TO47(-3320), .W62TO48(-1495), .W62TO49(11974), .W62TO50(15921), .W62TO51(-2291), .W62TO52(4092), .W62TO53(9714), .W62TO54(491), .W62TO55(22361), .W62TO56(-16067), .W62TO57(10326), .W62TO58(-5228), .W62TO59(7120), .W62TO60(11256), .W62TO61(-13918), .W62TO62(-14468), .W62TO63(-2574), .W62TO64(-18323), .W62TO65(1701), .W62TO66(7237), .W62TO67(21174), .W62TO68(-13038), .W62TO69(6813), .W62TO70(21495), .W62TO71(10475), .W62TO72(6763), .W62TO73(-4685), .W62TO74(-17908), .W62TO75(-4071), .W62TO76(21262), .W62TO77(-18113), .W62TO78(9423), .W62TO79(-9217), .W62TO80(6373), .W62TO81(-8384), .W62TO82(20774), .W62TO83(-11120), .W62TO84(4172), .W62TO85(2404), .W62TO86(-4444), .W62TO87(-11381), .W62TO88(13465), .W62TO89(-11665), .W62TO90(-10454), .W62TO91(-13810), .W62TO92(-9452), .W62TO93(9566), .W62TO94(13339), .W62TO95(-2319), .W62TO96(-11843), .W62TO97(-2226), .W62TO98(9651), .W62TO99(4904), .W63TO0(-2626), .W63TO1(-12820), .W63TO2(21694), .W63TO3(2428), .W63TO4(-3054), .W63TO5(-18219), .W63TO6(1672), .W63TO7(1433), .W63TO8(13374), .W63TO9(18731), .W63TO10(9780), .W63TO11(-8169), .W63TO12(-13830), .W63TO13(13939), .W63TO14(-14720), .W63TO15(-8705), .W63TO16(-18372), .W63TO17(-6407), .W63TO18(-9681), .W63TO19(7013), .W63TO20(16185), .W63TO21(-7526), .W63TO22(-7309), .W63TO23(-1703), .W63TO24(223), .W63TO25(3490), .W63TO26(12744), .W63TO27(325), .W63TO28(10483), .W63TO29(-14401), .W63TO30(7299), .W63TO31(-12219), .W63TO32(-10222), .W63TO33(-5007), .W63TO34(-7152), .W63TO35(4930), .W63TO36(-13189), .W63TO37(-14999), .W63TO38(-7893), .W63TO39(1986), .W63TO40(-14007), .W63TO41(2762), .W63TO42(14344), .W63TO43(13517), .W63TO44(-16847), .W63TO45(15097), .W63TO46(3235), .W63TO47(10202), .W63TO48(-8589), .W63TO49(-12150), .W63TO50(18851), .W63TO51(1010), .W63TO52(-14499), .W63TO53(1760), .W63TO54(-13952), .W63TO55(-10422), .W63TO56(16964), .W63TO57(14001), .W63TO58(12372), .W63TO59(14599), .W63TO60(14366), .W63TO61(-14626), .W63TO62(5335), .W63TO63(9120), .W63TO64(-6238), .W63TO65(-12340), .W63TO66(-5186), .W63TO67(8306), .W63TO68(14009), .W63TO69(6512), .W63TO70(9906), .W63TO71(8775), .W63TO72(13739), .W63TO73(8987), .W63TO74(15716), .W63TO75(-13906), .W63TO76(-15424), .W63TO77(-16030), .W63TO78(14032), .W63TO79(5038), .W63TO80(-2754), .W63TO81(-15342), .W63TO82(5781), .W63TO83(-4640), .W63TO84(3814), .W63TO85(-11150), .W63TO86(-12809), .W63TO87(-7512), .W63TO88(522), .W63TO89(-16395), .W63TO90(246), .W63TO91(-18269), .W63TO92(11550), .W63TO93(-16696), .W63TO94(7094), .W63TO95(-5076), .W63TO96(-8934), .W63TO97(-12630), .W63TO98(-8454), .W63TO99(-460)) layer0(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out0(con0[0]), .out1(con0[1]), .out2(con0[2]), .out3(con0[3]), .out4(con0[4]), .out5(con0[5]), .out6(con0[6]), .out7(con0[7]), .out8(con0[8]), .out9(con0[9]), .out10(con0[10]), .out11(con0[11]), .out12(con0[12]), .out13(con0[13]), .out14(con0[14]), .out15(con0[15]), .out16(con0[16]), .out17(con0[17]), .out18(con0[18]), .out19(con0[19]), .out20(con0[20]), .out21(con0[21]), .out22(con0[22]), .out23(con0[23]), .out24(con0[24]), .out25(con0[25]), .out26(con0[26]), .out27(con0[27]), .out28(con0[28]), .out29(con0[29]), .out30(con0[30]), .out31(con0[31]), .out32(con0[32]), .out33(con0[33]), .out34(con0[34]), .out35(con0[35]), .out36(con0[36]), .out37(con0[37]), .out38(con0[38]), .out39(con0[39]), .out40(con0[40]), .out41(con0[41]), .out42(con0[42]), .out43(con0[43]), .out44(con0[44]), .out45(con0[45]), .out46(con0[46]), .out47(con0[47]), .out48(con0[48]), .out49(con0[49]), .out50(con0[50]), .out51(con0[51]), .out52(con0[52]), .out53(con0[53]), .out54(con0[54]), .out55(con0[55]), .out56(con0[56]), .out57(con0[57]), .out58(con0[58]), .out59(con0[59]), .out60(con0[60]), .out61(con0[61]), .out62(con0[62]), .out63(con0[63]), .out64(con0[64]), .out65(con0[65]), .out66(con0[66]), .out67(con0[67]), .out68(con0[68]), .out69(con0[69]), .out70(con0[70]), .out71(con0[71]), .out72(con0[72]), .out73(con0[73]), .out74(con0[74]), .out75(con0[75]), .out76(con0[76]), .out77(con0[77]), .out78(con0[78]), .out79(con0[79]), .out80(con0[80]), .out81(con0[81]), .out82(con0[82]), .out83(con0[83]), .out84(con0[84]), .out85(con0[85]), .out86(con0[86]), .out87(con0[87]), .out88(con0[88]), .out89(con0[89]), .out90(con0[90]), .out91(con0[91]), .out92(con0[92]), .out93(con0[93]), .out94(con0[94]), .out95(con0[95]), .out96(con0[96]), .out97(con0[97]), .out98(con0[98]), .out99(con0[99]));
layer100in10out #(.W0TO0(26173), .W0TO1(21412), .W0TO2(25682), .W0TO3(26334), .W0TO4(6609), .W0TO5(-7002), .W0TO6(11470), .W0TO7(-14260), .W0TO8(29908), .W0TO9(6962), .W1TO0(-11349), .W1TO1(-14806), .W1TO2(-682), .W1TO3(6045), .W1TO4(-14691), .W1TO5(-3044), .W1TO6(-17890), .W1TO7(-8522), .W1TO8(12006), .W1TO9(-12549), .W2TO0(37785), .W2TO1(8063), .W2TO2(30081), .W2TO3(-12778), .W2TO4(-20582), .W2TO5(-6865), .W2TO6(-4027), .W2TO7(-7218), .W2TO8(531), .W2TO9(-12162), .W3TO0(-16729), .W3TO1(9444), .W3TO2(1688), .W3TO3(16710), .W3TO4(14224), .W3TO5(8021), .W3TO6(22730), .W3TO7(5014), .W3TO8(-2198), .W3TO9(19566), .W4TO0(17069), .W4TO1(17893), .W4TO2(30099), .W4TO3(-17001), .W4TO4(-2757), .W4TO5(-21845), .W4TO6(35920), .W4TO7(-10329), .W4TO8(-9496), .W4TO9(17618), .W5TO0(1142), .W5TO1(-16391), .W5TO2(735), .W5TO3(-1618), .W5TO4(11395), .W5TO5(46946), .W5TO6(-6950), .W5TO7(-14734), .W5TO8(-7381), .W5TO9(-22306), .W6TO0(-8104), .W6TO1(-27715), .W6TO2(-14207), .W6TO3(-2465), .W6TO4(-15527), .W6TO5(-21814), .W6TO6(-14897), .W6TO7(-16452), .W6TO8(15919), .W6TO9(4287), .W7TO0(15055), .W7TO1(-4847), .W7TO2(-1807), .W7TO3(11224), .W7TO4(-26416), .W7TO5(4734), .W7TO6(-10084), .W7TO7(51494), .W7TO8(-23348), .W7TO9(571), .W8TO0(-5813), .W8TO1(-15309), .W8TO2(-9022), .W8TO3(-23049), .W8TO4(8196), .W8TO5(-2857), .W8TO6(2635), .W8TO7(-2113), .W8TO8(32454), .W8TO9(-8208), .W9TO0(10452), .W9TO1(-21485), .W9TO2(16284), .W9TO3(-15175), .W9TO4(-25252), .W9TO5(-15573), .W9TO6(-11732), .W9TO7(-18537), .W9TO8(4449), .W9TO9(17628), .W10TO0(-7435), .W10TO1(1261), .W10TO2(11700), .W10TO3(-7210), .W10TO4(-17380), .W10TO5(1954), .W10TO6(7975), .W10TO7(15303), .W10TO8(-22469), .W10TO9(-26493), .W11TO0(-13224), .W11TO1(11084), .W11TO2(-7783), .W11TO3(-8090), .W11TO4(-21026), .W11TO5(-1023), .W11TO6(901), .W11TO7(-10686), .W11TO8(-11890), .W11TO9(8794), .W12TO0(-11477), .W12TO1(5946), .W12TO2(-13998), .W12TO3(15618), .W12TO4(13555), .W12TO5(-12684), .W12TO6(-36755), .W12TO7(16598), .W12TO8(16618), .W12TO9(-16422), .W13TO0(8773), .W13TO1(13033), .W13TO2(19365), .W13TO3(-8755), .W13TO4(-29915), .W13TO5(-26006), .W13TO6(-16144), .W13TO7(20253), .W13TO8(12900), .W13TO9(-13962), .W14TO0(-11022), .W14TO1(-13752), .W14TO2(-360), .W14TO3(3114), .W14TO4(6203), .W14TO5(10030), .W14TO6(-19047), .W14TO7(9454), .W14TO8(-17928), .W14TO9(181), .W15TO0(2286), .W15TO1(-24729), .W15TO2(12947), .W15TO3(3640), .W15TO4(-12648), .W15TO5(-27355), .W15TO6(-10071), .W15TO7(-8851), .W15TO8(15508), .W15TO9(19555), .W16TO0(-1873), .W16TO1(-15970), .W16TO2(-26504), .W16TO3(-24530), .W16TO4(14288), .W16TO5(17404), .W16TO6(4053), .W16TO7(7254), .W16TO8(-7847), .W16TO9(7071), .W17TO0(-23863), .W17TO1(36175), .W17TO2(3942), .W17TO3(134), .W17TO4(3859), .W17TO5(-7365), .W17TO6(-31682), .W17TO7(20414), .W17TO8(17236), .W17TO9(-24140), .W18TO0(-30742), .W18TO1(-3847), .W18TO2(1532), .W18TO3(8499), .W18TO4(-9433), .W18TO5(24382), .W18TO6(-2642), .W18TO7(-17426), .W18TO8(-13768), .W18TO9(9466), .W19TO0(-10982), .W19TO1(-2152), .W19TO2(29960), .W19TO3(40398), .W19TO4(-23587), .W19TO5(-24396), .W19TO6(-14179), .W19TO7(-18564), .W19TO8(5488), .W19TO9(-3768), .W20TO0(13148), .W20TO1(-5779), .W20TO2(-11242), .W20TO3(-17476), .W20TO4(17908), .W20TO5(21440), .W20TO6(-16858), .W20TO7(6658), .W20TO8(22691), .W20TO9(-22829), .W21TO0(-2441), .W21TO1(5563), .W21TO2(3192), .W21TO3(-16474), .W21TO4(-18743), .W21TO5(7556), .W21TO6(25041), .W21TO7(12897), .W21TO8(4948), .W21TO9(-14134), .W22TO0(8287), .W22TO1(24236), .W22TO2(15404), .W22TO3(2847), .W22TO4(-17526), .W22TO5(-21477), .W22TO6(11248), .W22TO7(-22361), .W22TO8(4524), .W22TO9(20580), .W23TO0(28048), .W23TO1(-3993), .W23TO2(7775), .W23TO3(19843), .W23TO4(-17817), .W23TO5(22453), .W23TO6(-4495), .W23TO7(-5083), .W23TO8(22878), .W23TO9(5952), .W24TO0(-15281), .W24TO1(-19703), .W24TO2(22519), .W24TO3(7893), .W24TO4(-24695), .W24TO5(-14978), .W24TO6(-15788), .W24TO7(19115), .W24TO8(15346), .W24TO9(16985), .W25TO0(-3547), .W25TO1(22920), .W25TO2(1233), .W25TO3(14974), .W25TO4(15958), .W25TO5(7678), .W25TO6(6188), .W25TO7(-2741), .W25TO8(-16952), .W25TO9(-1100), .W26TO0(19995), .W26TO1(5773), .W26TO2(-15620), .W26TO3(17410), .W26TO4(-10883), .W26TO5(-3032), .W26TO6(-1895), .W26TO7(11516), .W26TO8(-3433), .W26TO9(21933), .W27TO0(22686), .W27TO1(895), .W27TO2(-3093), .W27TO3(6585), .W27TO4(1330), .W27TO5(-6665), .W27TO6(3913), .W27TO7(14733), .W27TO8(27473), .W27TO9(23038), .W28TO0(-12081), .W28TO1(-5312), .W28TO2(7800), .W28TO3(6066), .W28TO4(-16976), .W28TO5(-9547), .W28TO6(-7329), .W28TO7(22703), .W28TO8(16156), .W28TO9(16548), .W29TO0(26639), .W29TO1(-44798), .W29TO2(-769), .W29TO3(-13317), .W29TO4(36182), .W29TO5(-7259), .W29TO6(-17653), .W29TO7(32119), .W29TO8(3820), .W29TO9(29194), .W30TO0(13595), .W30TO1(-11959), .W30TO2(-9188), .W30TO3(-7299), .W30TO4(-1857), .W30TO5(-21016), .W30TO6(34422), .W30TO7(-6348), .W30TO8(25401), .W30TO9(1549), .W31TO0(-15095), .W31TO1(-5408), .W31TO2(-12972), .W31TO3(-10367), .W31TO4(28604), .W31TO5(-15725), .W31TO6(11442), .W31TO7(-3046), .W31TO8(18126), .W31TO9(-29712), .W32TO0(-2591), .W32TO1(-16072), .W32TO2(-18345), .W32TO3(-13039), .W32TO4(16020), .W32TO5(-23661), .W32TO6(12675), .W32TO7(-11278), .W32TO8(-29109), .W32TO9(-15644), .W33TO0(9295), .W33TO1(-19504), .W33TO2(-28634), .W33TO3(14202), .W33TO4(9667), .W33TO5(26451), .W33TO6(23023), .W33TO7(12652), .W33TO8(20200), .W33TO9(-18743), .W34TO0(-8995), .W34TO1(6855), .W34TO2(-13567), .W34TO3(-6517), .W34TO4(-807), .W34TO5(21484), .W34TO6(5101), .W34TO7(-13142), .W34TO8(6345), .W34TO9(18185), .W35TO0(8700), .W35TO1(1129), .W35TO2(-13024), .W35TO3(-20069), .W35TO4(-21057), .W35TO5(4184), .W35TO6(-382), .W35TO7(-19065), .W35TO8(89), .W35TO9(17869), .W36TO0(3), .W36TO1(5587), .W36TO2(10903), .W36TO3(-37360), .W36TO4(13609), .W36TO5(26975), .W36TO6(11670), .W36TO7(-21415), .W36TO8(15848), .W36TO9(-13645), .W37TO0(-8890), .W37TO1(13750), .W37TO2(-9187), .W37TO3(-8106), .W37TO4(-26027), .W37TO5(12112), .W37TO6(-21390), .W37TO7(-21709), .W37TO8(-12624), .W37TO9(1268), .W38TO0(-4013), .W38TO1(-16944), .W38TO2(-10794), .W38TO3(3056), .W38TO4(4025), .W38TO5(-22824), .W38TO6(7751), .W38TO7(-2771), .W38TO8(-20819), .W38TO9(-24730), .W39TO0(-7012), .W39TO1(-15309), .W39TO2(3718), .W39TO3(16285), .W39TO4(28819), .W39TO5(-16638), .W39TO6(-1447), .W39TO7(3197), .W39TO8(-15295), .W39TO9(13624), .W40TO0(-16802), .W40TO1(9607), .W40TO2(24246), .W40TO3(24492), .W40TO4(6987), .W40TO5(15829), .W40TO6(23825), .W40TO7(-9267), .W40TO8(26072), .W40TO9(16083), .W41TO0(37359), .W41TO1(-30697), .W41TO2(13965), .W41TO3(-8780), .W41TO4(-11186), .W41TO5(-21110), .W41TO6(7226), .W41TO7(-21841), .W41TO8(24974), .W41TO9(-25661), .W42TO0(10050), .W42TO1(23186), .W42TO2(3173), .W42TO3(22362), .W42TO4(1389), .W42TO5(17086), .W42TO6(-12350), .W42TO7(26470), .W42TO8(21512), .W42TO9(18349), .W43TO0(-707), .W43TO1(16711), .W43TO2(7205), .W43TO3(13104), .W43TO4(3270), .W43TO5(-11353), .W43TO6(-12382), .W43TO7(-30417), .W43TO8(5079), .W43TO9(-5243), .W44TO0(18249), .W44TO1(-9020), .W44TO2(11274), .W44TO3(6961), .W44TO4(-7882), .W44TO5(-22302), .W44TO6(-15320), .W44TO7(-6036), .W44TO8(-19290), .W44TO9(16536), .W45TO0(26227), .W45TO1(10169), .W45TO2(-13588), .W45TO3(-3042), .W45TO4(-17670), .W45TO5(11705), .W45TO6(21919), .W45TO7(24411), .W45TO8(11991), .W45TO9(-5083), .W46TO0(9794), .W46TO1(-25), .W46TO2(-3427), .W46TO3(27945), .W46TO4(19882), .W46TO5(22660), .W46TO6(-1073), .W46TO7(8349), .W46TO8(2918), .W46TO9(23505), .W47TO0(-21111), .W47TO1(4603), .W47TO2(5581), .W47TO3(20687), .W47TO4(-24282), .W47TO5(-21684), .W47TO6(-25348), .W47TO7(18978), .W47TO8(23674), .W47TO9(35947), .W48TO0(15126), .W48TO1(-13210), .W48TO2(2953), .W48TO3(20371), .W48TO4(7605), .W48TO5(-18042), .W48TO6(21641), .W48TO7(-1298), .W48TO8(-1173), .W48TO9(19126), .W49TO0(6755), .W49TO1(2744), .W49TO2(-44667), .W49TO3(18709), .W49TO4(-14366), .W49TO5(1554), .W49TO6(-8986), .W49TO7(-29224), .W49TO8(19924), .W49TO9(-11122), .W50TO0(-18513), .W50TO1(-12549), .W50TO2(10775), .W50TO3(5765), .W50TO4(4365), .W50TO5(-16305), .W50TO6(-7285), .W50TO7(-9944), .W50TO8(9694), .W50TO9(13518), .W51TO0(6899), .W51TO1(-29237), .W51TO2(-19217), .W51TO3(-6954), .W51TO4(15023), .W51TO5(-20243), .W51TO6(-4734), .W51TO7(15922), .W51TO8(10510), .W51TO9(8414), .W52TO0(-8770), .W52TO1(-32987), .W52TO2(16455), .W52TO3(-13025), .W52TO4(-24692), .W52TO5(20254), .W52TO6(13168), .W52TO7(-8215), .W52TO8(9565), .W52TO9(-1889), .W53TO0(-39661), .W53TO1(12917), .W53TO2(16863), .W53TO3(-8178), .W53TO4(-30569), .W53TO5(9624), .W53TO6(18555), .W53TO7(5459), .W53TO8(23125), .W53TO9(-21930), .W54TO0(4449), .W54TO1(-23072), .W54TO2(-25313), .W54TO3(-22132), .W54TO4(3131), .W54TO5(4202), .W54TO6(42833), .W54TO7(9452), .W54TO8(-7141), .W54TO9(5610), .W55TO0(-20803), .W55TO1(22040), .W55TO2(270), .W55TO3(-4868), .W55TO4(-5767), .W55TO5(-23527), .W55TO6(12931), .W55TO7(11529), .W55TO8(411), .W55TO9(7546), .W56TO0(-1448), .W56TO1(-13221), .W56TO2(-19294), .W56TO3(-9340), .W56TO4(-17064), .W56TO5(13831), .W56TO6(-10640), .W56TO7(16101), .W56TO8(-16441), .W56TO9(-7419), .W57TO0(22562), .W57TO1(17506), .W57TO2(16679), .W57TO3(-17020), .W57TO4(24958), .W57TO5(-14780), .W57TO6(5089), .W57TO7(-4112), .W57TO8(6215), .W57TO9(-974), .W58TO0(19244), .W58TO1(-4981), .W58TO2(35113), .W58TO3(-14103), .W58TO4(8692), .W58TO5(-4473), .W58TO6(-259), .W58TO7(15049), .W58TO8(18199), .W58TO9(15339), .W59TO0(31403), .W59TO1(-21808), .W59TO2(17004), .W59TO3(5177), .W59TO4(-9757), .W59TO5(-7366), .W59TO6(24091), .W59TO7(5357), .W59TO8(-32082), .W59TO9(-39202), .W60TO0(-21252), .W60TO1(49502), .W60TO2(-16001), .W60TO3(-26720), .W60TO4(26625), .W60TO5(-12075), .W60TO6(19994), .W60TO7(-10448), .W60TO8(-24875), .W60TO9(726), .W61TO0(7631), .W61TO1(11766), .W61TO2(-9160), .W61TO3(7516), .W61TO4(-16214), .W61TO5(-29978), .W61TO6(-7443), .W61TO7(39639), .W61TO8(22072), .W61TO9(11685), .W62TO0(-11923), .W62TO1(-18143), .W62TO2(6492), .W62TO3(-4458), .W62TO4(5707), .W62TO5(8446), .W62TO6(-12089), .W62TO7(24149), .W62TO8(27824), .W62TO9(21867), .W63TO0(22050), .W63TO1(-24114), .W63TO2(7799), .W63TO3(405), .W63TO4(-35229), .W63TO5(1935), .W63TO6(-4125), .W63TO7(-13534), .W63TO8(-15748), .W63TO9(-7520), .W64TO0(-1740), .W64TO1(-4692), .W64TO2(32056), .W64TO3(-17082), .W64TO4(-6428), .W64TO5(14579), .W64TO6(-11860), .W64TO7(-1938), .W64TO8(-4207), .W64TO9(-5846), .W65TO0(-19851), .W65TO1(20881), .W65TO2(13038), .W65TO3(-3913), .W65TO4(28973), .W65TO5(5143), .W65TO6(-17191), .W65TO7(-20434), .W65TO8(-16663), .W65TO9(-11973), .W66TO0(26019), .W66TO1(16069), .W66TO2(20912), .W66TO3(25887), .W66TO4(17946), .W66TO5(23953), .W66TO6(714), .W66TO7(2781), .W66TO8(-9095), .W66TO9(-3038), .W67TO0(-13979), .W67TO1(-10127), .W67TO2(33664), .W67TO3(23207), .W67TO4(-7644), .W67TO5(4475), .W67TO6(14466), .W67TO7(-10237), .W67TO8(-32348), .W67TO9(-22402), .W68TO0(-12117), .W68TO1(-10278), .W68TO2(-26474), .W68TO3(-20937), .W68TO4(-17956), .W68TO5(6929), .W68TO6(5812), .W68TO7(-24396), .W68TO8(-27089), .W68TO9(-20657), .W69TO0(-2268), .W69TO1(-12580), .W69TO2(15683), .W69TO3(14058), .W69TO4(10376), .W69TO5(7009), .W69TO6(-20711), .W69TO7(16246), .W69TO8(-20143), .W69TO9(-12513), .W70TO0(-12186), .W70TO1(-15791), .W70TO2(15432), .W70TO3(-9508), .W70TO4(-6798), .W70TO5(-27010), .W70TO6(27262), .W70TO7(-18172), .W70TO8(22855), .W70TO9(27471), .W71TO0(20701), .W71TO1(-7660), .W71TO2(-21674), .W71TO3(22387), .W71TO4(4378), .W71TO5(-5168), .W71TO6(-6235), .W71TO7(1377), .W71TO8(2657), .W71TO9(19349), .W72TO0(16369), .W72TO1(-8813), .W72TO2(-20292), .W72TO3(-13119), .W72TO4(-11696), .W72TO5(-11263), .W72TO6(-16392), .W72TO7(-27622), .W72TO8(-22737), .W72TO9(3382), .W73TO0(-17278), .W73TO1(12041), .W73TO2(21902), .W73TO3(-11695), .W73TO4(-12838), .W73TO5(16388), .W73TO6(-2665), .W73TO7(6673), .W73TO8(5660), .W73TO9(-13649), .W74TO0(-7726), .W74TO1(-1679), .W74TO2(20505), .W74TO3(22495), .W74TO4(26033), .W74TO5(18642), .W74TO6(-80), .W74TO7(22338), .W74TO8(-6572), .W74TO9(-1361), .W75TO0(7672), .W75TO1(5495), .W75TO2(-18667), .W75TO3(8958), .W75TO4(665), .W75TO5(22126), .W75TO6(13791), .W75TO7(-13572), .W75TO8(18283), .W75TO9(18281), .W76TO0(10043), .W76TO1(-7284), .W76TO2(12030), .W76TO3(20173), .W76TO4(-5459), .W76TO5(11266), .W76TO6(-3529), .W76TO7(-25651), .W76TO8(-6758), .W76TO9(-26619), .W77TO0(-934), .W77TO1(2390), .W77TO2(-7878), .W77TO3(-2127), .W77TO4(-2080), .W77TO5(24408), .W77TO6(-1407), .W77TO7(17742), .W77TO8(10444), .W77TO9(32), .W78TO0(2156), .W78TO1(12845), .W78TO2(20681), .W78TO3(-29567), .W78TO4(17045), .W78TO5(-22778), .W78TO6(-4469), .W78TO7(19568), .W78TO8(-34152), .W78TO9(-40187), .W79TO0(16904), .W79TO1(624), .W79TO2(-6096), .W79TO3(29153), .W79TO4(-2212), .W79TO5(6120), .W79TO6(1323), .W79TO7(2610), .W79TO8(-11173), .W79TO9(-25656), .W80TO0(20008), .W80TO1(5684), .W80TO2(14368), .W80TO3(-12596), .W80TO4(8405), .W80TO5(-23113), .W80TO6(8031), .W80TO7(-20896), .W80TO8(39619), .W80TO9(-16504), .W81TO0(3004), .W81TO1(-18553), .W81TO2(-15083), .W81TO3(-11597), .W81TO4(-25776), .W81TO5(365), .W81TO6(-7279), .W81TO7(-13179), .W81TO8(2479), .W81TO9(-21674), .W82TO0(-35395), .W82TO1(9791), .W82TO2(7889), .W82TO3(16513), .W82TO4(-32008), .W82TO5(18340), .W82TO6(26098), .W82TO7(-35882), .W82TO8(24922), .W82TO9(29281), .W83TO0(-2902), .W83TO1(-23407), .W83TO2(3803), .W83TO3(36248), .W83TO4(-8315), .W83TO5(16712), .W83TO6(-26453), .W83TO7(-4688), .W83TO8(-25955), .W83TO9(32075), .W84TO0(-17734), .W84TO1(35498), .W84TO2(-4089), .W84TO3(-36092), .W84TO4(21771), .W84TO5(-26765), .W84TO6(5213), .W84TO7(8839), .W84TO8(14440), .W84TO9(25041), .W85TO0(-17441), .W85TO1(12714), .W85TO2(-20592), .W85TO3(-7297), .W85TO4(-13165), .W85TO5(-22783), .W85TO6(-1190), .W85TO7(11264), .W85TO8(-22538), .W85TO9(8024), .W86TO0(2746), .W86TO1(23473), .W86TO2(-15263), .W86TO3(13257), .W86TO4(8068), .W86TO5(609), .W86TO6(-15069), .W86TO7(-5163), .W86TO8(-23187), .W86TO9(19921), .W87TO0(24863), .W87TO1(-22298), .W87TO2(-13658), .W87TO3(-15355), .W87TO4(14933), .W87TO5(22562), .W87TO6(2549), .W87TO7(-6305), .W87TO8(17100), .W87TO9(-4174), .W88TO0(-15389), .W88TO1(34711), .W88TO2(-23374), .W88TO3(3902), .W88TO4(-1305), .W88TO5(-16204), .W88TO6(19598), .W88TO7(397), .W88TO8(7676), .W88TO9(13519), .W89TO0(7222), .W89TO1(25017), .W89TO2(15980), .W89TO3(-11903), .W89TO4(-40884), .W89TO5(-12872), .W89TO6(16318), .W89TO7(-14268), .W89TO8(7700), .W89TO9(-18401), .W90TO0(-9655), .W90TO1(15945), .W90TO2(-4954), .W90TO3(-21701), .W90TO4(-6132), .W90TO5(-17097), .W90TO6(-24774), .W90TO7(-21264), .W90TO8(-11721), .W90TO9(-22623), .W91TO0(15426), .W91TO1(8074), .W91TO2(-2616), .W91TO3(40047), .W91TO4(-3755), .W91TO5(-22748), .W91TO6(-3250), .W91TO7(-15192), .W91TO8(-4429), .W91TO9(-12472), .W92TO0(-14263), .W92TO1(8482), .W92TO2(11529), .W92TO3(690), .W92TO4(9135), .W92TO5(4691), .W92TO6(5462), .W92TO7(14922), .W92TO8(12004), .W92TO9(-326), .W93TO0(-31992), .W93TO1(2075), .W93TO2(6051), .W93TO3(17613), .W93TO4(19160), .W93TO5(-12354), .W93TO6(14429), .W93TO7(24486), .W93TO8(21388), .W93TO9(-37841), .W94TO0(2053), .W94TO1(15255), .W94TO2(21080), .W94TO3(12912), .W94TO4(18717), .W94TO5(-16571), .W94TO6(23509), .W94TO7(25272), .W94TO8(2373), .W94TO9(10299), .W95TO0(-21915), .W95TO1(8347), .W95TO2(9396), .W95TO3(24519), .W95TO4(12352), .W95TO5(-24165), .W95TO6(7946), .W95TO7(2073), .W95TO8(220), .W95TO9(-33821), .W96TO0(-11920), .W96TO1(-2957), .W96TO2(16225), .W96TO3(-3432), .W96TO4(-1390), .W96TO5(4862), .W96TO6(-23360), .W96TO7(3372), .W96TO8(14123), .W96TO9(-12176), .W97TO0(23159), .W97TO1(-5143), .W97TO2(185), .W97TO3(-1902), .W97TO4(-17414), .W97TO5(-3806), .W97TO6(-2989), .W97TO7(6584), .W97TO8(-7983), .W97TO9(-10641), .W98TO0(-2688), .W98TO1(798), .W98TO2(15542), .W98TO3(-14506), .W98TO4(14723), .W98TO5(-26488), .W98TO6(2465), .W98TO7(-34254), .W98TO8(9184), .W98TO9(8903), .W99TO0(-17988), .W99TO1(-28038), .W99TO2(-26118), .W99TO3(-13254), .W99TO4(8546), .W99TO5(145), .W99TO6(-6541), .W99TO7(143), .W99TO8(14059), .W99TO9(-19670)) layer1(.clk(clk), .rst(rst), .in0(con0[0]), .in1(con0[1]), .in2(con0[2]), .in3(con0[3]), .in4(con0[4]), .in5(con0[5]), .in6(con0[6]), .in7(con0[7]), .in8(con0[8]), .in9(con0[9]), .in10(con0[10]), .in11(con0[11]), .in12(con0[12]), .in13(con0[13]), .in14(con0[14]), .in15(con0[15]), .in16(con0[16]), .in17(con0[17]), .in18(con0[18]), .in19(con0[19]), .in20(con0[20]), .in21(con0[21]), .in22(con0[22]), .in23(con0[23]), .in24(con0[24]), .in25(con0[25]), .in26(con0[26]), .in27(con0[27]), .in28(con0[28]), .in29(con0[29]), .in30(con0[30]), .in31(con0[31]), .in32(con0[32]), .in33(con0[33]), .in34(con0[34]), .in35(con0[35]), .in36(con0[36]), .in37(con0[37]), .in38(con0[38]), .in39(con0[39]), .in40(con0[40]), .in41(con0[41]), .in42(con0[42]), .in43(con0[43]), .in44(con0[44]), .in45(con0[45]), .in46(con0[46]), .in47(con0[47]), .in48(con0[48]), .in49(con0[49]), .in50(con0[50]), .in51(con0[51]), .in52(con0[52]), .in53(con0[53]), .in54(con0[54]), .in55(con0[55]), .in56(con0[56]), .in57(con0[57]), .in58(con0[58]), .in59(con0[59]), .in60(con0[60]), .in61(con0[61]), .in62(con0[62]), .in63(con0[63]), .in64(con0[64]), .in65(con0[65]), .in66(con0[66]), .in67(con0[67]), .in68(con0[68]), .in69(con0[69]), .in70(con0[70]), .in71(con0[71]), .in72(con0[72]), .in73(con0[73]), .in74(con0[74]), .in75(con0[75]), .in76(con0[76]), .in77(con0[77]), .in78(con0[78]), .in79(con0[79]), .in80(con0[80]), .in81(con0[81]), .in82(con0[82]), .in83(con0[83]), .in84(con0[84]), .in85(con0[85]), .in86(con0[86]), .in87(con0[87]), .in88(con0[88]), .in89(con0[89]), .in90(con0[90]), .in91(con0[91]), .in92(con0[92]), .in93(con0[93]), .in94(con0[94]), .in95(con0[95]), .in96(con0[96]), .in97(con0[97]), .in98(con0[98]), .in99(con0[99]), .out0(out0), .out1(out1), .out2(out2), .out3(out3), .out4(out4), .out5(out5), .out6(out6), .out7(out7), .out8(out8), .out9(out9));

endmodule

module testbench_digits;

logic clk;
logic rst;

reg [15:0] net_in0, net_in1, net_in2, net_in3, net_in4, net_in5, net_in6, net_in7, net_in8, net_in9, net_in10, net_in11, net_in12, net_in13, net_in14, net_in15, net_in16, net_in17, net_in18, net_in19, net_in20, net_in21, net_in22, net_in23, net_in24, net_in25, net_in26, net_in27, net_in28, net_in29, net_in30, net_in31, net_in32, net_in33, net_in34, net_in35, net_in36, net_in37, net_in38, net_in39, net_in40, net_in41, net_in42, net_in43, net_in44, net_in45, net_in46, net_in47, net_in48, net_in49, net_in50, net_in51, net_in52, net_in53, net_in54, net_in55, net_in56, net_in57, net_in58, net_in59, net_in60, net_in61, net_in62, net_in63;
wire [15:0] net_out0, net_out1, net_out2, net_out3, net_out4, net_out5, net_out6, net_out7, net_out8, net_out9;

network net(.clk(clk), .rst(rst), .in0(net_in0), .in1(net_in1), .in2(net_in2), .in3(net_in3), .in4(net_in4), .in5(net_in5), .in6(net_in6), .in7(net_in7), .in8(net_in8), .in9(net_in9), .in10(net_in10), .in11(net_in11), .in12(net_in12), .in13(net_in13), .in14(net_in14), .in15(net_in15), .in16(net_in16), .in17(net_in17), .in18(net_in18), .in19(net_in19), .in20(net_in20), .in21(net_in21), .in22(net_in22), .in23(net_in23), .in24(net_in24), .in25(net_in25), .in26(net_in26), .in27(net_in27), .in28(net_in28), .in29(net_in29), .in30(net_in30), .in31(net_in31), .in32(net_in32), .in33(net_in33), .in34(net_in34), .in35(net_in35), .in36(net_in36), .in37(net_in37), .in38(net_in38), .in39(net_in39), .in40(net_in40), .in41(net_in41), .in42(net_in42), .in43(net_in43), .in44(net_in44), .in45(net_in45), .in46(net_in46), .in47(net_in47), .in48(net_in48), .in49(net_in49), .in50(net_in50), .in51(net_in51), .in52(net_in52), .in53(net_in53), .in54(net_in54), .in55(net_in55), .in56(net_in56), .in57(net_in57), .in58(net_in58), .in59(net_in59), .in60(net_in60), .in61(net_in61), .in62(net_in62), .in63(net_in63), .out0(net_out0), .out1(net_out1), .out2(net_out2), .out3(net_out3), .out4(net_out4), .out5(net_out5), .out6(net_out6), .out7(net_out7), .out8(net_out8), .out9(net_out9));

task test;
input [15:0] in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63;
begin
    net_in0 = in0;
    net_in1 = in1;
    net_in2 = in2;
    net_in3 = in3;
    net_in4 = in4;
    net_in5 = in5;
    net_in6 = in6;
    net_in7 = in7;
    net_in8 = in8;
    net_in9 = in9;
    net_in10 = in10;
    net_in11 = in11;
    net_in12 = in12;
    net_in13 = in13;
    net_in14 = in14;
    net_in15 = in15;
    net_in16 = in16;
    net_in17 = in17;
    net_in18 = in18;
    net_in19 = in19;
    net_in20 = in20;
    net_in21 = in21;
    net_in22 = in22;
    net_in23 = in23;
    net_in24 = in24;
    net_in25 = in25;
    net_in26 = in26;
    net_in27 = in27;
    net_in28 = in28;
    net_in29 = in29;
    net_in30 = in30;
    net_in31 = in31;
    net_in32 = in32;
    net_in33 = in33;
    net_in34 = in34;
    net_in35 = in35;
    net_in36 = in36;
    net_in37 = in37;
    net_in38 = in38;
    net_in39 = in39;
    net_in40 = in40;
    net_in41 = in41;
    net_in42 = in42;
    net_in43 = in43;
    net_in44 = in44;
    net_in45 = in45;
    net_in46 = in46;
    net_in47 = in47;
    net_in48 = in48;
    net_in49 = in49;
    net_in50 = in50;
    net_in51 = in51;
    net_in52 = in52;
    net_in53 = in53;
    net_in54 = in54;
    net_in55 = in55;
    net_in56 = in56;
    net_in57 = in57;
    net_in58 = in58;
    net_in59 = in59;
    net_in60 = in60;
    net_in61 = in61;
    net_in62 = in62;
    net_in63 = in63;
    #10000000

    $write("%d ", net_out0);
    $write("%d ", net_out1);
    $write("%d ", net_out2);
    $write("%d ", net_out3);
    $write("%d ", net_out4);
    $write("%d ", net_out5);
    $write("%d ", net_out6);
    $write("%d ", net_out7);
    $write("%d ", net_out8);
    $write("%d ", net_out9);
    $display();
end
endtask

initial begin
    test(0, 0, 1, 15, 15, 2, 0, 0, 0, 0, 3, 12, 16, 6, 0, 0, 0, 0, 0, 4, 16, 4, 0, 0, 0, 0, 3, 8, 16, 4, 0, 0, 0, 10, 16, 16, 16, 16, 8, 0, 0, 8, 11, 14, 14, 5, 1, 0, 0, 0, 0, 15, 6, 0, 0, 0, 0, 0, 1, 15, 2, 0, 0, 0);
    test(0, 0, 13, 13, 8, 2, 0, 0, 0, 5, 16, 16, 16, 12, 0, 0, 0, 1, 15, 12, 0, 0, 0, 0, 0, 0, 12, 13, 7, 1, 0, 0, 0, 0, 8, 16, 16, 12, 0, 0, 0, 0, 0, 4, 9, 16, 3, 0, 0, 0, 1, 5, 14, 15, 1, 0, 0, 0, 10, 16, 16, 6, 0, 0);
    test(0, 0, 14, 12, 12, 12, 6, 0, 0, 2, 15, 8, 8, 8, 4, 0, 0, 5, 12, 0, 0, 0, 0, 0, 0, 8, 16, 12, 11, 7, 0, 0, 0, 1, 4, 4, 9, 15, 7, 0, 0, 0, 0, 0, 0, 8, 8, 0, 0, 1, 11, 4, 5, 14, 7, 0, 0, 0, 12, 16, 16, 8, 1, 0);
    test(0, 0, 0, 5, 13, 16, 8, 0, 0, 0, 8, 15, 6, 7, 14, 0, 0, 2, 16, 1, 1, 11, 10, 0, 0, 4, 16, 15, 16, 16, 6, 0, 0, 0, 4, 4, 5, 15, 1, 0, 0, 0, 0, 0, 9, 8, 0, 0, 0, 0, 0, 2, 15, 1, 0, 0, 0, 0, 0, 6, 10, 0, 0, 0);
    test(0, 0, 5, 13, 16, 14, 0, 0, 0, 1, 14, 8, 5, 16, 2, 0, 0, 0, 1, 0, 2, 15, 2, 0, 0, 0, 0, 2, 8, 15, 3, 0, 0, 0, 0, 15, 16, 13, 8, 0, 0, 0, 0, 6, 14, 0, 0, 0, 0, 0, 0, 13, 7, 0, 0, 0, 0, 0, 7, 14, 0, 0, 0, 0);
    test(0, 2, 13, 16, 16, 16, 15, 2, 0, 8, 16, 12, 8, 4, 1, 0, 0, 5, 16, 13, 1, 0, 0, 0, 0, 0, 8, 16, 8, 0, 0, 0, 0, 0, 0, 10, 16, 0, 0, 0, 0, 0, 0, 9, 16, 0, 0, 0, 0, 0, 3, 13, 12, 0, 0, 0, 0, 2, 16, 16, 6, 0, 0, 0);
    test(0, 1, 12, 15, 16, 13, 1, 0, 0, 4, 16, 15, 7, 15, 4, 0, 0, 0, 16, 6, 11, 15, 2, 0, 0, 0, 9, 16, 15, 4, 0, 0, 0, 0, 8, 16, 8, 0, 0, 0, 0, 0, 15, 15, 11, 0, 0, 0, 0, 2, 16, 10, 12, 0, 0, 0, 0, 2, 13, 16, 10, 0, 0, 0);
    test(0, 3, 12, 12, 14, 4, 0, 0, 0, 1, 13, 4, 4, 0, 0, 0, 0, 4, 14, 4, 3, 0, 0, 0, 0, 5, 13, 12, 14, 10, 0, 0, 0, 0, 0, 0, 0, 11, 6, 0, 0, 0, 0, 0, 0, 4, 8, 0, 0, 0, 6, 2, 0, 8, 8, 0, 0, 2, 13, 16, 16, 16, 2, 0);
    test(0, 0, 4, 14, 16, 5, 0, 0, 0, 4, 16, 16, 16, 8, 0, 0, 0, 12, 12, 0, 15, 8, 0, 0, 0, 2, 1, 5, 16, 13, 1, 0, 0, 0, 0, 1, 11, 15, 11, 0, 0, 0, 0, 0, 0, 11, 12, 0, 0, 0, 2, 13, 12, 16, 7, 0, 0, 0, 3, 16, 15, 8, 0, 0);
    test(0, 0, 5, 8, 11, 5, 0, 0, 0, 0, 13, 16, 12, 12, 0, 0, 0, 1, 16, 9, 0, 9, 3, 0, 0, 3, 16, 6, 0, 6, 6, 0, 0, 3, 11, 1, 0, 5, 6, 0, 0, 0, 12, 0, 0, 11, 6, 0, 0, 0, 14, 5, 12, 15, 1, 0, 0, 0, 6, 16, 13, 2, 0, 0);
end
endmodule
