module neuron65in(clk, rst, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, out);

parameter signed BIAS = 0;
parameter signed W0 = 0;
parameter signed W1 = 0;
parameter signed W2 = 0;
parameter signed W3 = 0;
parameter signed W4 = 0;
parameter signed W5 = 0;
parameter signed W6 = 0;
parameter signed W7 = 0;
parameter signed W8 = 0;
parameter signed W9 = 0;
parameter signed W10 = 0;
parameter signed W11 = 0;
parameter signed W12 = 0;
parameter signed W13 = 0;
parameter signed W14 = 0;
parameter signed W15 = 0;
parameter signed W16 = 0;
parameter signed W17 = 0;
parameter signed W18 = 0;
parameter signed W19 = 0;
parameter signed W20 = 0;
parameter signed W21 = 0;
parameter signed W22 = 0;
parameter signed W23 = 0;
parameter signed W24 = 0;
parameter signed W25 = 0;
parameter signed W26 = 0;
parameter signed W27 = 0;
parameter signed W28 = 0;
parameter signed W29 = 0;
parameter signed W30 = 0;
parameter signed W31 = 0;
parameter signed W32 = 0;
parameter signed W33 = 0;
parameter signed W34 = 0;
parameter signed W35 = 0;
parameter signed W36 = 0;
parameter signed W37 = 0;
parameter signed W38 = 0;
parameter signed W39 = 0;
parameter signed W40 = 0;
parameter signed W41 = 0;
parameter signed W42 = 0;
parameter signed W43 = 0;
parameter signed W44 = 0;
parameter signed W45 = 0;
parameter signed W46 = 0;
parameter signed W47 = 0;
parameter signed W48 = 0;
parameter signed W49 = 0;
parameter signed W50 = 0;
parameter signed W51 = 0;
parameter signed W52 = 0;
parameter signed W53 = 0;
parameter signed W54 = 0;
parameter signed W55 = 0;
parameter signed W56 = 0;
parameter signed W57 = 0;
parameter signed W58 = 0;
parameter signed W59 = 0;
parameter signed W60 = 0;
parameter signed W61 = 0;
parameter signed W62 = 0;
parameter signed W63 = 0;
parameter signed W64 = 0;

input wire clk;
input wire rst;

input signed [15:0] in0;
input signed [15:0] in1;
input signed [15:0] in2;
input signed [15:0] in3;
input signed [15:0] in4;
input signed [15:0] in5;
input signed [15:0] in6;
input signed [15:0] in7;
input signed [15:0] in8;
input signed [15:0] in9;
input signed [15:0] in10;
input signed [15:0] in11;
input signed [15:0] in12;
input signed [15:0] in13;
input signed [15:0] in14;
input signed [15:0] in15;
input signed [15:0] in16;
input signed [15:0] in17;
input signed [15:0] in18;
input signed [15:0] in19;
input signed [15:0] in20;
input signed [15:0] in21;
input signed [15:0] in22;
input signed [15:0] in23;
input signed [15:0] in24;
input signed [15:0] in25;
input signed [15:0] in26;
input signed [15:0] in27;
input signed [15:0] in28;
input signed [15:0] in29;
input signed [15:0] in30;
input signed [15:0] in31;
input signed [15:0] in32;
input signed [15:0] in33;
input signed [15:0] in34;
input signed [15:0] in35;
input signed [15:0] in36;
input signed [15:0] in37;
input signed [15:0] in38;
input signed [15:0] in39;
input signed [15:0] in40;
input signed [15:0] in41;
input signed [15:0] in42;
input signed [15:0] in43;
input signed [15:0] in44;
input signed [15:0] in45;
input signed [15:0] in46;
input signed [15:0] in47;
input signed [15:0] in48;
input signed [15:0] in49;
input signed [15:0] in50;
input signed [15:0] in51;
input signed [15:0] in52;
input signed [15:0] in53;
input signed [15:0] in54;
input signed [15:0] in55;
input signed [15:0] in56;
input signed [15:0] in57;
input signed [15:0] in58;
input signed [15:0] in59;
input signed [15:0] in60;
input signed [15:0] in61;
input signed [15:0] in62;
input signed [15:0] in63;
input signed [15:0] in64;

output reg signed [15:0] out;

reg signed [31:0] x;
reg signed [31:0] abs_x;
reg signed [31:0] y;
reg signed [31:0] sum_0_0;
reg signed [31:0] sum_0_1;
reg signed [31:0] sum_0_2;
reg signed [31:0] sum_0_3;
reg signed [31:0] sum_0_4;
reg signed [31:0] sum_0_5;
reg signed [31:0] sum_0_6;
reg signed [31:0] sum_0_7;
reg signed [31:0] sum_0_8;
reg signed [31:0] sum_0_9;
reg signed [31:0] sum_0_10;
reg signed [31:0] sum_0_11;
reg signed [31:0] sum_0_12;
reg signed [31:0] sum_0_13;
reg signed [31:0] sum_0_14;
reg signed [31:0] sum_0_15;
reg signed [31:0] sum_0_16;
reg signed [31:0] sum_0_17;
reg signed [31:0] sum_0_18;
reg signed [31:0] sum_0_19;
reg signed [31:0] sum_0_20;
reg signed [31:0] sum_0_21;
reg signed [31:0] sum_0_22;
reg signed [31:0] sum_0_23;
reg signed [31:0] sum_0_24;
reg signed [31:0] sum_0_25;
reg signed [31:0] sum_0_26;
reg signed [31:0] sum_0_27;
reg signed [31:0] sum_0_28;
reg signed [31:0] sum_0_29;
reg signed [31:0] sum_0_30;
reg signed [31:0] sum_0_31;
reg signed [31:0] sum_0_32;
reg signed [31:0] sum_1_0;
reg signed [31:0] sum_1_1;
reg signed [31:0] sum_1_2;
reg signed [31:0] sum_1_3;
reg signed [31:0] sum_1_4;
reg signed [31:0] sum_1_5;
reg signed [31:0] sum_1_6;
reg signed [31:0] sum_1_7;
reg signed [31:0] sum_1_8;
reg signed [31:0] sum_1_9;
reg signed [31:0] sum_1_10;
reg signed [31:0] sum_1_11;
reg signed [31:0] sum_1_12;
reg signed [31:0] sum_1_13;
reg signed [31:0] sum_1_14;
reg signed [31:0] sum_1_15;
reg signed [31:0] sum_2_0;
reg signed [31:0] sum_2_1;
reg signed [31:0] sum_2_2;
reg signed [31:0] sum_2_3;
reg signed [31:0] sum_2_4;
reg signed [31:0] sum_2_5;
reg signed [31:0] sum_2_6;
reg signed [31:0] sum_2_7;
reg signed [31:0] sum_3_0;
reg signed [31:0] sum_3_1;
reg signed [31:0] sum_3_2;
reg signed [31:0] sum_3_3;
reg signed [31:0] sum_4_0;
reg signed [31:0] sum_4_1;
reg signed [31:0] sum_5_0;
always @* begin
    sum_0_0 <= (in0 * W0 + 500) / 1000 + (in1 * W1 + 500) / 1000;
    sum_0_1 <= (in2 * W2 + 500) / 1000 + (in3 * W3 + 500) / 1000;
    sum_0_2 <= (in4 * W4 + 500) / 1000 + (in5 * W5 + 500) / 1000;
    sum_0_3 <= (in6 * W6 + 500) / 1000 + (in7 * W7 + 500) / 1000;
    sum_0_4 <= (in8 * W8 + 500) / 1000 + (in9 * W9 + 500) / 1000;
    sum_0_5 <= (in10 * W10 + 500) / 1000 + (in11 * W11 + 500) / 1000;
    sum_0_6 <= (in12 * W12 + 500) / 1000 + (in13 * W13 + 500) / 1000;
    sum_0_7 <= (in14 * W14 + 500) / 1000 + (in15 * W15 + 500) / 1000;
    sum_0_8 <= (in16 * W16 + 500) / 1000 + (in17 * W17 + 500) / 1000;
    sum_0_9 <= (in18 * W18 + 500) / 1000 + (in19 * W19 + 500) / 1000;
    sum_0_10 <= (in20 * W20 + 500) / 1000 + (in21 * W21 + 500) / 1000;
    sum_0_11 <= (in22 * W22 + 500) / 1000 + (in23 * W23 + 500) / 1000;
    sum_0_12 <= (in24 * W24 + 500) / 1000 + (in25 * W25 + 500) / 1000;
    sum_0_13 <= (in26 * W26 + 500) / 1000 + (in27 * W27 + 500) / 1000;
    sum_0_14 <= (in28 * W28 + 500) / 1000 + (in29 * W29 + 500) / 1000;
    sum_0_15 <= (in30 * W30 + 500) / 1000 + (in31 * W31 + 500) / 1000;
    sum_0_16 <= (in32 * W32 + 500) / 1000 + (in33 * W33 + 500) / 1000;
    sum_0_17 <= (in34 * W34 + 500) / 1000 + (in35 * W35 + 500) / 1000;
    sum_0_18 <= (in36 * W36 + 500) / 1000 + (in37 * W37 + 500) / 1000;
    sum_0_19 <= (in38 * W38 + 500) / 1000 + (in39 * W39 + 500) / 1000;
    sum_0_20 <= (in40 * W40 + 500) / 1000 + (in41 * W41 + 500) / 1000;
    sum_0_21 <= (in42 * W42 + 500) / 1000 + (in43 * W43 + 500) / 1000;
    sum_0_22 <= (in44 * W44 + 500) / 1000 + (in45 * W45 + 500) / 1000;
    sum_0_23 <= (in46 * W46 + 500) / 1000 + (in47 * W47 + 500) / 1000;
    sum_0_24 <= (in48 * W48 + 500) / 1000 + (in49 * W49 + 500) / 1000;
    sum_0_25 <= (in50 * W50 + 500) / 1000 + (in51 * W51 + 500) / 1000;
    sum_0_26 <= (in52 * W52 + 500) / 1000 + (in53 * W53 + 500) / 1000;
    sum_0_27 <= (in54 * W54 + 500) / 1000 + (in55 * W55 + 500) / 1000;
    sum_0_28 <= (in56 * W56 + 500) / 1000 + (in57 * W57 + 500) / 1000;
    sum_0_29 <= (in58 * W58 + 500) / 1000 + (in59 * W59 + 500) / 1000;
    sum_0_30 <= (in60 * W60 + 500) / 1000 + (in61 * W61 + 500) / 1000;
    sum_0_31 <= (in62 * W62 + 500) / 1000 + (in63 * W63 + 500) / 1000;
    sum_0_32 <= (in64 * W64 + 500) / 1000 + BIAS;
    sum_1_0 <= sum_0_0 + sum_0_1;
    sum_1_1 <= sum_0_2 + sum_0_3;
    sum_1_2 <= sum_0_4 + sum_0_5;
    sum_1_3 <= sum_0_6 + sum_0_7;
    sum_1_4 <= sum_0_8 + sum_0_9;
    sum_1_5 <= sum_0_10 + sum_0_11;
    sum_1_6 <= sum_0_12 + sum_0_13;
    sum_1_7 <= sum_0_14 + sum_0_15;
    sum_1_8 <= sum_0_16 + sum_0_17;
    sum_1_9 <= sum_0_18 + sum_0_19;
    sum_1_10 <= sum_0_20 + sum_0_21;
    sum_1_11 <= sum_0_22 + sum_0_23;
    sum_1_12 <= sum_0_24 + sum_0_25;
    sum_1_13 <= sum_0_26 + sum_0_27;
    sum_1_14 <= sum_0_28 + sum_0_29;
    sum_1_15 <= sum_0_30 + sum_0_31 + sum_0_32;
    sum_2_0 <= sum_1_0 + sum_1_1;
    sum_2_1 <= sum_1_2 + sum_1_3;
    sum_2_2 <= sum_1_4 + sum_1_5;
    sum_2_3 <= sum_1_6 + sum_1_7;
    sum_2_4 <= sum_1_8 + sum_1_9;
    sum_2_5 <= sum_1_10 + sum_1_11;
    sum_2_6 <= sum_1_12 + sum_1_13;
    sum_2_7 <= sum_1_14 + sum_1_15;
    sum_3_0 <= sum_2_0 + sum_2_1;
    sum_3_1 <= sum_2_2 + sum_2_3;
    sum_3_2 <= sum_2_4 + sum_2_5;
    sum_3_3 <= sum_2_6 + sum_2_7;
    sum_4_0 <= sum_3_0 + sum_3_1;
    sum_4_1 <= sum_3_2 + sum_3_3;
    sum_5_0 <= sum_4_0 + sum_4_1;
    x <= sum_5_0;
    abs_x = x < 0 ? -x : x;
    if (abs_x >= 5000) y = 1000;
    else if (abs_x >= 2375) y = 31 * abs_x / 1000 + 844;
    else if (abs_x >= 1000) y = 125 * abs_x / 1000 + 625;
    else y = 250 * abs_x / 1000 + 500;
    out = x < 0 ? 1000 - y : y;
end

endmodule

module neuron64in(clk, rst, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, out);

parameter signed BIAS = 0;
parameter signed W0 = 0;
parameter signed W1 = 0;
parameter signed W2 = 0;
parameter signed W3 = 0;
parameter signed W4 = 0;
parameter signed W5 = 0;
parameter signed W6 = 0;
parameter signed W7 = 0;
parameter signed W8 = 0;
parameter signed W9 = 0;
parameter signed W10 = 0;
parameter signed W11 = 0;
parameter signed W12 = 0;
parameter signed W13 = 0;
parameter signed W14 = 0;
parameter signed W15 = 0;
parameter signed W16 = 0;
parameter signed W17 = 0;
parameter signed W18 = 0;
parameter signed W19 = 0;
parameter signed W20 = 0;
parameter signed W21 = 0;
parameter signed W22 = 0;
parameter signed W23 = 0;
parameter signed W24 = 0;
parameter signed W25 = 0;
parameter signed W26 = 0;
parameter signed W27 = 0;
parameter signed W28 = 0;
parameter signed W29 = 0;
parameter signed W30 = 0;
parameter signed W31 = 0;
parameter signed W32 = 0;
parameter signed W33 = 0;
parameter signed W34 = 0;
parameter signed W35 = 0;
parameter signed W36 = 0;
parameter signed W37 = 0;
parameter signed W38 = 0;
parameter signed W39 = 0;
parameter signed W40 = 0;
parameter signed W41 = 0;
parameter signed W42 = 0;
parameter signed W43 = 0;
parameter signed W44 = 0;
parameter signed W45 = 0;
parameter signed W46 = 0;
parameter signed W47 = 0;
parameter signed W48 = 0;
parameter signed W49 = 0;
parameter signed W50 = 0;
parameter signed W51 = 0;
parameter signed W52 = 0;
parameter signed W53 = 0;
parameter signed W54 = 0;
parameter signed W55 = 0;
parameter signed W56 = 0;
parameter signed W57 = 0;
parameter signed W58 = 0;
parameter signed W59 = 0;
parameter signed W60 = 0;
parameter signed W61 = 0;
parameter signed W62 = 0;
parameter signed W63 = 0;

input wire clk;
input wire rst;

input signed [15:0] in0;
input signed [15:0] in1;
input signed [15:0] in2;
input signed [15:0] in3;
input signed [15:0] in4;
input signed [15:0] in5;
input signed [15:0] in6;
input signed [15:0] in7;
input signed [15:0] in8;
input signed [15:0] in9;
input signed [15:0] in10;
input signed [15:0] in11;
input signed [15:0] in12;
input signed [15:0] in13;
input signed [15:0] in14;
input signed [15:0] in15;
input signed [15:0] in16;
input signed [15:0] in17;
input signed [15:0] in18;
input signed [15:0] in19;
input signed [15:0] in20;
input signed [15:0] in21;
input signed [15:0] in22;
input signed [15:0] in23;
input signed [15:0] in24;
input signed [15:0] in25;
input signed [15:0] in26;
input signed [15:0] in27;
input signed [15:0] in28;
input signed [15:0] in29;
input signed [15:0] in30;
input signed [15:0] in31;
input signed [15:0] in32;
input signed [15:0] in33;
input signed [15:0] in34;
input signed [15:0] in35;
input signed [15:0] in36;
input signed [15:0] in37;
input signed [15:0] in38;
input signed [15:0] in39;
input signed [15:0] in40;
input signed [15:0] in41;
input signed [15:0] in42;
input signed [15:0] in43;
input signed [15:0] in44;
input signed [15:0] in45;
input signed [15:0] in46;
input signed [15:0] in47;
input signed [15:0] in48;
input signed [15:0] in49;
input signed [15:0] in50;
input signed [15:0] in51;
input signed [15:0] in52;
input signed [15:0] in53;
input signed [15:0] in54;
input signed [15:0] in55;
input signed [15:0] in56;
input signed [15:0] in57;
input signed [15:0] in58;
input signed [15:0] in59;
input signed [15:0] in60;
input signed [15:0] in61;
input signed [15:0] in62;
input signed [15:0] in63;

output reg signed [15:0] out;

reg signed [31:0] x;
reg signed [31:0] abs_x;
reg signed [31:0] y;
reg signed [31:0] sum_0_0;
reg signed [31:0] sum_0_1;
reg signed [31:0] sum_0_2;
reg signed [31:0] sum_0_3;
reg signed [31:0] sum_0_4;
reg signed [31:0] sum_0_5;
reg signed [31:0] sum_0_6;
reg signed [31:0] sum_0_7;
reg signed [31:0] sum_0_8;
reg signed [31:0] sum_0_9;
reg signed [31:0] sum_0_10;
reg signed [31:0] sum_0_11;
reg signed [31:0] sum_0_12;
reg signed [31:0] sum_0_13;
reg signed [31:0] sum_0_14;
reg signed [31:0] sum_0_15;
reg signed [31:0] sum_0_16;
reg signed [31:0] sum_0_17;
reg signed [31:0] sum_0_18;
reg signed [31:0] sum_0_19;
reg signed [31:0] sum_0_20;
reg signed [31:0] sum_0_21;
reg signed [31:0] sum_0_22;
reg signed [31:0] sum_0_23;
reg signed [31:0] sum_0_24;
reg signed [31:0] sum_0_25;
reg signed [31:0] sum_0_26;
reg signed [31:0] sum_0_27;
reg signed [31:0] sum_0_28;
reg signed [31:0] sum_0_29;
reg signed [31:0] sum_0_30;
reg signed [31:0] sum_0_31;
reg signed [31:0] sum_1_0;
reg signed [31:0] sum_1_1;
reg signed [31:0] sum_1_2;
reg signed [31:0] sum_1_3;
reg signed [31:0] sum_1_4;
reg signed [31:0] sum_1_5;
reg signed [31:0] sum_1_6;
reg signed [31:0] sum_1_7;
reg signed [31:0] sum_1_8;
reg signed [31:0] sum_1_9;
reg signed [31:0] sum_1_10;
reg signed [31:0] sum_1_11;
reg signed [31:0] sum_1_12;
reg signed [31:0] sum_1_13;
reg signed [31:0] sum_1_14;
reg signed [31:0] sum_1_15;
reg signed [31:0] sum_2_0;
reg signed [31:0] sum_2_1;
reg signed [31:0] sum_2_2;
reg signed [31:0] sum_2_3;
reg signed [31:0] sum_2_4;
reg signed [31:0] sum_2_5;
reg signed [31:0] sum_2_6;
reg signed [31:0] sum_2_7;
reg signed [31:0] sum_3_0;
reg signed [31:0] sum_3_1;
reg signed [31:0] sum_3_2;
reg signed [31:0] sum_3_3;
reg signed [31:0] sum_4_0;
reg signed [31:0] sum_4_1;
reg signed [31:0] sum_5_0;
always @* begin
    sum_0_0 <= (in0 * W0 + 500) / 1000 + (in1 * W1 + 500) / 1000;
    sum_0_1 <= (in2 * W2 + 500) / 1000 + (in3 * W3 + 500) / 1000;
    sum_0_2 <= (in4 * W4 + 500) / 1000 + (in5 * W5 + 500) / 1000;
    sum_0_3 <= (in6 * W6 + 500) / 1000 + (in7 * W7 + 500) / 1000;
    sum_0_4 <= (in8 * W8 + 500) / 1000 + (in9 * W9 + 500) / 1000;
    sum_0_5 <= (in10 * W10 + 500) / 1000 + (in11 * W11 + 500) / 1000;
    sum_0_6 <= (in12 * W12 + 500) / 1000 + (in13 * W13 + 500) / 1000;
    sum_0_7 <= (in14 * W14 + 500) / 1000 + (in15 * W15 + 500) / 1000;
    sum_0_8 <= (in16 * W16 + 500) / 1000 + (in17 * W17 + 500) / 1000;
    sum_0_9 <= (in18 * W18 + 500) / 1000 + (in19 * W19 + 500) / 1000;
    sum_0_10 <= (in20 * W20 + 500) / 1000 + (in21 * W21 + 500) / 1000;
    sum_0_11 <= (in22 * W22 + 500) / 1000 + (in23 * W23 + 500) / 1000;
    sum_0_12 <= (in24 * W24 + 500) / 1000 + (in25 * W25 + 500) / 1000;
    sum_0_13 <= (in26 * W26 + 500) / 1000 + (in27 * W27 + 500) / 1000;
    sum_0_14 <= (in28 * W28 + 500) / 1000 + (in29 * W29 + 500) / 1000;
    sum_0_15 <= (in30 * W30 + 500) / 1000 + (in31 * W31 + 500) / 1000;
    sum_0_16 <= (in32 * W32 + 500) / 1000 + (in33 * W33 + 500) / 1000;
    sum_0_17 <= (in34 * W34 + 500) / 1000 + (in35 * W35 + 500) / 1000;
    sum_0_18 <= (in36 * W36 + 500) / 1000 + (in37 * W37 + 500) / 1000;
    sum_0_19 <= (in38 * W38 + 500) / 1000 + (in39 * W39 + 500) / 1000;
    sum_0_20 <= (in40 * W40 + 500) / 1000 + (in41 * W41 + 500) / 1000;
    sum_0_21 <= (in42 * W42 + 500) / 1000 + (in43 * W43 + 500) / 1000;
    sum_0_22 <= (in44 * W44 + 500) / 1000 + (in45 * W45 + 500) / 1000;
    sum_0_23 <= (in46 * W46 + 500) / 1000 + (in47 * W47 + 500) / 1000;
    sum_0_24 <= (in48 * W48 + 500) / 1000 + (in49 * W49 + 500) / 1000;
    sum_0_25 <= (in50 * W50 + 500) / 1000 + (in51 * W51 + 500) / 1000;
    sum_0_26 <= (in52 * W52 + 500) / 1000 + (in53 * W53 + 500) / 1000;
    sum_0_27 <= (in54 * W54 + 500) / 1000 + (in55 * W55 + 500) / 1000;
    sum_0_28 <= (in56 * W56 + 500) / 1000 + (in57 * W57 + 500) / 1000;
    sum_0_29 <= (in58 * W58 + 500) / 1000 + (in59 * W59 + 500) / 1000;
    sum_0_30 <= (in60 * W60 + 500) / 1000 + (in61 * W61 + 500) / 1000;
    sum_0_31 <= (in62 * W62 + 500) / 1000 + (in63 * W63 + 500) / 1000 + BIAS;
    sum_1_0 <= sum_0_0 + sum_0_1;
    sum_1_1 <= sum_0_2 + sum_0_3;
    sum_1_2 <= sum_0_4 + sum_0_5;
    sum_1_3 <= sum_0_6 + sum_0_7;
    sum_1_4 <= sum_0_8 + sum_0_9;
    sum_1_5 <= sum_0_10 + sum_0_11;
    sum_1_6 <= sum_0_12 + sum_0_13;
    sum_1_7 <= sum_0_14 + sum_0_15;
    sum_1_8 <= sum_0_16 + sum_0_17;
    sum_1_9 <= sum_0_18 + sum_0_19;
    sum_1_10 <= sum_0_20 + sum_0_21;
    sum_1_11 <= sum_0_22 + sum_0_23;
    sum_1_12 <= sum_0_24 + sum_0_25;
    sum_1_13 <= sum_0_26 + sum_0_27;
    sum_1_14 <= sum_0_28 + sum_0_29;
    sum_1_15 <= sum_0_30 + sum_0_31;
    sum_2_0 <= sum_1_0 + sum_1_1;
    sum_2_1 <= sum_1_2 + sum_1_3;
    sum_2_2 <= sum_1_4 + sum_1_5;
    sum_2_3 <= sum_1_6 + sum_1_7;
    sum_2_4 <= sum_1_8 + sum_1_9;
    sum_2_5 <= sum_1_10 + sum_1_11;
    sum_2_6 <= sum_1_12 + sum_1_13;
    sum_2_7 <= sum_1_14 + sum_1_15;
    sum_3_0 <= sum_2_0 + sum_2_1;
    sum_3_1 <= sum_2_2 + sum_2_3;
    sum_3_2 <= sum_2_4 + sum_2_5;
    sum_3_3 <= sum_2_6 + sum_2_7;
    sum_4_0 <= sum_3_0 + sum_3_1;
    sum_4_1 <= sum_3_2 + sum_3_3;
    sum_5_0 <= sum_4_0 + sum_4_1;
    x <= sum_5_0;
    abs_x = x < 0 ? -x : x;
    if (abs_x >= 5000) y = 1000;
    else if (abs_x >= 2375) y = 31 * abs_x / 1000 + 844;
    else if (abs_x >= 1000) y = 125 * abs_x / 1000 + 625;
    else y = 250 * abs_x / 1000 + 500;
    out = x < 0 ? 1000 - y : y;
end

endmodule

module layer65in64out(clk, rst, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, out0, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13, out14, out15, out16, out17, out18, out19, out20, out21, out22, out23, out24, out25, out26, out27, out28, out29, out30, out31, out32, out33, out34, out35, out36, out37, out38, out39, out40, out41, out42, out43, out44, out45, out46, out47, out48, out49, out50, out51, out52, out53, out54, out55, out56, out57, out58, out59, out60, out61, out62, out63);

parameter signed BIAS0 = 0;
parameter signed BIAS1 = 0;
parameter signed BIAS2 = 0;
parameter signed BIAS3 = 0;
parameter signed BIAS4 = 0;
parameter signed BIAS5 = 0;
parameter signed BIAS6 = 0;
parameter signed BIAS7 = 0;
parameter signed BIAS8 = 0;
parameter signed BIAS9 = 0;
parameter signed BIAS10 = 0;
parameter signed BIAS11 = 0;
parameter signed BIAS12 = 0;
parameter signed BIAS13 = 0;
parameter signed BIAS14 = 0;
parameter signed BIAS15 = 0;
parameter signed BIAS16 = 0;
parameter signed BIAS17 = 0;
parameter signed BIAS18 = 0;
parameter signed BIAS19 = 0;
parameter signed BIAS20 = 0;
parameter signed BIAS21 = 0;
parameter signed BIAS22 = 0;
parameter signed BIAS23 = 0;
parameter signed BIAS24 = 0;
parameter signed BIAS25 = 0;
parameter signed BIAS26 = 0;
parameter signed BIAS27 = 0;
parameter signed BIAS28 = 0;
parameter signed BIAS29 = 0;
parameter signed BIAS30 = 0;
parameter signed BIAS31 = 0;
parameter signed BIAS32 = 0;
parameter signed BIAS33 = 0;
parameter signed BIAS34 = 0;
parameter signed BIAS35 = 0;
parameter signed BIAS36 = 0;
parameter signed BIAS37 = 0;
parameter signed BIAS38 = 0;
parameter signed BIAS39 = 0;
parameter signed BIAS40 = 0;
parameter signed BIAS41 = 0;
parameter signed BIAS42 = 0;
parameter signed BIAS43 = 0;
parameter signed BIAS44 = 0;
parameter signed BIAS45 = 0;
parameter signed BIAS46 = 0;
parameter signed BIAS47 = 0;
parameter signed BIAS48 = 0;
parameter signed BIAS49 = 0;
parameter signed BIAS50 = 0;
parameter signed BIAS51 = 0;
parameter signed BIAS52 = 0;
parameter signed BIAS53 = 0;
parameter signed BIAS54 = 0;
parameter signed BIAS55 = 0;
parameter signed BIAS56 = 0;
parameter signed BIAS57 = 0;
parameter signed BIAS58 = 0;
parameter signed BIAS59 = 0;
parameter signed BIAS60 = 0;
parameter signed BIAS61 = 0;
parameter signed BIAS62 = 0;
parameter signed BIAS63 = 0;
parameter signed W0TO0 = 0;
parameter signed W0TO1 = 0;
parameter signed W0TO2 = 0;
parameter signed W0TO3 = 0;
parameter signed W0TO4 = 0;
parameter signed W0TO5 = 0;
parameter signed W0TO6 = 0;
parameter signed W0TO7 = 0;
parameter signed W0TO8 = 0;
parameter signed W0TO9 = 0;
parameter signed W0TO10 = 0;
parameter signed W0TO11 = 0;
parameter signed W0TO12 = 0;
parameter signed W0TO13 = 0;
parameter signed W0TO14 = 0;
parameter signed W0TO15 = 0;
parameter signed W0TO16 = 0;
parameter signed W0TO17 = 0;
parameter signed W0TO18 = 0;
parameter signed W0TO19 = 0;
parameter signed W0TO20 = 0;
parameter signed W0TO21 = 0;
parameter signed W0TO22 = 0;
parameter signed W0TO23 = 0;
parameter signed W0TO24 = 0;
parameter signed W0TO25 = 0;
parameter signed W0TO26 = 0;
parameter signed W0TO27 = 0;
parameter signed W0TO28 = 0;
parameter signed W0TO29 = 0;
parameter signed W0TO30 = 0;
parameter signed W0TO31 = 0;
parameter signed W0TO32 = 0;
parameter signed W0TO33 = 0;
parameter signed W0TO34 = 0;
parameter signed W0TO35 = 0;
parameter signed W0TO36 = 0;
parameter signed W0TO37 = 0;
parameter signed W0TO38 = 0;
parameter signed W0TO39 = 0;
parameter signed W0TO40 = 0;
parameter signed W0TO41 = 0;
parameter signed W0TO42 = 0;
parameter signed W0TO43 = 0;
parameter signed W0TO44 = 0;
parameter signed W0TO45 = 0;
parameter signed W0TO46 = 0;
parameter signed W0TO47 = 0;
parameter signed W0TO48 = 0;
parameter signed W0TO49 = 0;
parameter signed W0TO50 = 0;
parameter signed W0TO51 = 0;
parameter signed W0TO52 = 0;
parameter signed W0TO53 = 0;
parameter signed W0TO54 = 0;
parameter signed W0TO55 = 0;
parameter signed W0TO56 = 0;
parameter signed W0TO57 = 0;
parameter signed W0TO58 = 0;
parameter signed W0TO59 = 0;
parameter signed W0TO60 = 0;
parameter signed W0TO61 = 0;
parameter signed W0TO62 = 0;
parameter signed W0TO63 = 0;
parameter signed W1TO0 = 0;
parameter signed W1TO1 = 0;
parameter signed W1TO2 = 0;
parameter signed W1TO3 = 0;
parameter signed W1TO4 = 0;
parameter signed W1TO5 = 0;
parameter signed W1TO6 = 0;
parameter signed W1TO7 = 0;
parameter signed W1TO8 = 0;
parameter signed W1TO9 = 0;
parameter signed W1TO10 = 0;
parameter signed W1TO11 = 0;
parameter signed W1TO12 = 0;
parameter signed W1TO13 = 0;
parameter signed W1TO14 = 0;
parameter signed W1TO15 = 0;
parameter signed W1TO16 = 0;
parameter signed W1TO17 = 0;
parameter signed W1TO18 = 0;
parameter signed W1TO19 = 0;
parameter signed W1TO20 = 0;
parameter signed W1TO21 = 0;
parameter signed W1TO22 = 0;
parameter signed W1TO23 = 0;
parameter signed W1TO24 = 0;
parameter signed W1TO25 = 0;
parameter signed W1TO26 = 0;
parameter signed W1TO27 = 0;
parameter signed W1TO28 = 0;
parameter signed W1TO29 = 0;
parameter signed W1TO30 = 0;
parameter signed W1TO31 = 0;
parameter signed W1TO32 = 0;
parameter signed W1TO33 = 0;
parameter signed W1TO34 = 0;
parameter signed W1TO35 = 0;
parameter signed W1TO36 = 0;
parameter signed W1TO37 = 0;
parameter signed W1TO38 = 0;
parameter signed W1TO39 = 0;
parameter signed W1TO40 = 0;
parameter signed W1TO41 = 0;
parameter signed W1TO42 = 0;
parameter signed W1TO43 = 0;
parameter signed W1TO44 = 0;
parameter signed W1TO45 = 0;
parameter signed W1TO46 = 0;
parameter signed W1TO47 = 0;
parameter signed W1TO48 = 0;
parameter signed W1TO49 = 0;
parameter signed W1TO50 = 0;
parameter signed W1TO51 = 0;
parameter signed W1TO52 = 0;
parameter signed W1TO53 = 0;
parameter signed W1TO54 = 0;
parameter signed W1TO55 = 0;
parameter signed W1TO56 = 0;
parameter signed W1TO57 = 0;
parameter signed W1TO58 = 0;
parameter signed W1TO59 = 0;
parameter signed W1TO60 = 0;
parameter signed W1TO61 = 0;
parameter signed W1TO62 = 0;
parameter signed W1TO63 = 0;
parameter signed W2TO0 = 0;
parameter signed W2TO1 = 0;
parameter signed W2TO2 = 0;
parameter signed W2TO3 = 0;
parameter signed W2TO4 = 0;
parameter signed W2TO5 = 0;
parameter signed W2TO6 = 0;
parameter signed W2TO7 = 0;
parameter signed W2TO8 = 0;
parameter signed W2TO9 = 0;
parameter signed W2TO10 = 0;
parameter signed W2TO11 = 0;
parameter signed W2TO12 = 0;
parameter signed W2TO13 = 0;
parameter signed W2TO14 = 0;
parameter signed W2TO15 = 0;
parameter signed W2TO16 = 0;
parameter signed W2TO17 = 0;
parameter signed W2TO18 = 0;
parameter signed W2TO19 = 0;
parameter signed W2TO20 = 0;
parameter signed W2TO21 = 0;
parameter signed W2TO22 = 0;
parameter signed W2TO23 = 0;
parameter signed W2TO24 = 0;
parameter signed W2TO25 = 0;
parameter signed W2TO26 = 0;
parameter signed W2TO27 = 0;
parameter signed W2TO28 = 0;
parameter signed W2TO29 = 0;
parameter signed W2TO30 = 0;
parameter signed W2TO31 = 0;
parameter signed W2TO32 = 0;
parameter signed W2TO33 = 0;
parameter signed W2TO34 = 0;
parameter signed W2TO35 = 0;
parameter signed W2TO36 = 0;
parameter signed W2TO37 = 0;
parameter signed W2TO38 = 0;
parameter signed W2TO39 = 0;
parameter signed W2TO40 = 0;
parameter signed W2TO41 = 0;
parameter signed W2TO42 = 0;
parameter signed W2TO43 = 0;
parameter signed W2TO44 = 0;
parameter signed W2TO45 = 0;
parameter signed W2TO46 = 0;
parameter signed W2TO47 = 0;
parameter signed W2TO48 = 0;
parameter signed W2TO49 = 0;
parameter signed W2TO50 = 0;
parameter signed W2TO51 = 0;
parameter signed W2TO52 = 0;
parameter signed W2TO53 = 0;
parameter signed W2TO54 = 0;
parameter signed W2TO55 = 0;
parameter signed W2TO56 = 0;
parameter signed W2TO57 = 0;
parameter signed W2TO58 = 0;
parameter signed W2TO59 = 0;
parameter signed W2TO60 = 0;
parameter signed W2TO61 = 0;
parameter signed W2TO62 = 0;
parameter signed W2TO63 = 0;
parameter signed W3TO0 = 0;
parameter signed W3TO1 = 0;
parameter signed W3TO2 = 0;
parameter signed W3TO3 = 0;
parameter signed W3TO4 = 0;
parameter signed W3TO5 = 0;
parameter signed W3TO6 = 0;
parameter signed W3TO7 = 0;
parameter signed W3TO8 = 0;
parameter signed W3TO9 = 0;
parameter signed W3TO10 = 0;
parameter signed W3TO11 = 0;
parameter signed W3TO12 = 0;
parameter signed W3TO13 = 0;
parameter signed W3TO14 = 0;
parameter signed W3TO15 = 0;
parameter signed W3TO16 = 0;
parameter signed W3TO17 = 0;
parameter signed W3TO18 = 0;
parameter signed W3TO19 = 0;
parameter signed W3TO20 = 0;
parameter signed W3TO21 = 0;
parameter signed W3TO22 = 0;
parameter signed W3TO23 = 0;
parameter signed W3TO24 = 0;
parameter signed W3TO25 = 0;
parameter signed W3TO26 = 0;
parameter signed W3TO27 = 0;
parameter signed W3TO28 = 0;
parameter signed W3TO29 = 0;
parameter signed W3TO30 = 0;
parameter signed W3TO31 = 0;
parameter signed W3TO32 = 0;
parameter signed W3TO33 = 0;
parameter signed W3TO34 = 0;
parameter signed W3TO35 = 0;
parameter signed W3TO36 = 0;
parameter signed W3TO37 = 0;
parameter signed W3TO38 = 0;
parameter signed W3TO39 = 0;
parameter signed W3TO40 = 0;
parameter signed W3TO41 = 0;
parameter signed W3TO42 = 0;
parameter signed W3TO43 = 0;
parameter signed W3TO44 = 0;
parameter signed W3TO45 = 0;
parameter signed W3TO46 = 0;
parameter signed W3TO47 = 0;
parameter signed W3TO48 = 0;
parameter signed W3TO49 = 0;
parameter signed W3TO50 = 0;
parameter signed W3TO51 = 0;
parameter signed W3TO52 = 0;
parameter signed W3TO53 = 0;
parameter signed W3TO54 = 0;
parameter signed W3TO55 = 0;
parameter signed W3TO56 = 0;
parameter signed W3TO57 = 0;
parameter signed W3TO58 = 0;
parameter signed W3TO59 = 0;
parameter signed W3TO60 = 0;
parameter signed W3TO61 = 0;
parameter signed W3TO62 = 0;
parameter signed W3TO63 = 0;
parameter signed W4TO0 = 0;
parameter signed W4TO1 = 0;
parameter signed W4TO2 = 0;
parameter signed W4TO3 = 0;
parameter signed W4TO4 = 0;
parameter signed W4TO5 = 0;
parameter signed W4TO6 = 0;
parameter signed W4TO7 = 0;
parameter signed W4TO8 = 0;
parameter signed W4TO9 = 0;
parameter signed W4TO10 = 0;
parameter signed W4TO11 = 0;
parameter signed W4TO12 = 0;
parameter signed W4TO13 = 0;
parameter signed W4TO14 = 0;
parameter signed W4TO15 = 0;
parameter signed W4TO16 = 0;
parameter signed W4TO17 = 0;
parameter signed W4TO18 = 0;
parameter signed W4TO19 = 0;
parameter signed W4TO20 = 0;
parameter signed W4TO21 = 0;
parameter signed W4TO22 = 0;
parameter signed W4TO23 = 0;
parameter signed W4TO24 = 0;
parameter signed W4TO25 = 0;
parameter signed W4TO26 = 0;
parameter signed W4TO27 = 0;
parameter signed W4TO28 = 0;
parameter signed W4TO29 = 0;
parameter signed W4TO30 = 0;
parameter signed W4TO31 = 0;
parameter signed W4TO32 = 0;
parameter signed W4TO33 = 0;
parameter signed W4TO34 = 0;
parameter signed W4TO35 = 0;
parameter signed W4TO36 = 0;
parameter signed W4TO37 = 0;
parameter signed W4TO38 = 0;
parameter signed W4TO39 = 0;
parameter signed W4TO40 = 0;
parameter signed W4TO41 = 0;
parameter signed W4TO42 = 0;
parameter signed W4TO43 = 0;
parameter signed W4TO44 = 0;
parameter signed W4TO45 = 0;
parameter signed W4TO46 = 0;
parameter signed W4TO47 = 0;
parameter signed W4TO48 = 0;
parameter signed W4TO49 = 0;
parameter signed W4TO50 = 0;
parameter signed W4TO51 = 0;
parameter signed W4TO52 = 0;
parameter signed W4TO53 = 0;
parameter signed W4TO54 = 0;
parameter signed W4TO55 = 0;
parameter signed W4TO56 = 0;
parameter signed W4TO57 = 0;
parameter signed W4TO58 = 0;
parameter signed W4TO59 = 0;
parameter signed W4TO60 = 0;
parameter signed W4TO61 = 0;
parameter signed W4TO62 = 0;
parameter signed W4TO63 = 0;
parameter signed W5TO0 = 0;
parameter signed W5TO1 = 0;
parameter signed W5TO2 = 0;
parameter signed W5TO3 = 0;
parameter signed W5TO4 = 0;
parameter signed W5TO5 = 0;
parameter signed W5TO6 = 0;
parameter signed W5TO7 = 0;
parameter signed W5TO8 = 0;
parameter signed W5TO9 = 0;
parameter signed W5TO10 = 0;
parameter signed W5TO11 = 0;
parameter signed W5TO12 = 0;
parameter signed W5TO13 = 0;
parameter signed W5TO14 = 0;
parameter signed W5TO15 = 0;
parameter signed W5TO16 = 0;
parameter signed W5TO17 = 0;
parameter signed W5TO18 = 0;
parameter signed W5TO19 = 0;
parameter signed W5TO20 = 0;
parameter signed W5TO21 = 0;
parameter signed W5TO22 = 0;
parameter signed W5TO23 = 0;
parameter signed W5TO24 = 0;
parameter signed W5TO25 = 0;
parameter signed W5TO26 = 0;
parameter signed W5TO27 = 0;
parameter signed W5TO28 = 0;
parameter signed W5TO29 = 0;
parameter signed W5TO30 = 0;
parameter signed W5TO31 = 0;
parameter signed W5TO32 = 0;
parameter signed W5TO33 = 0;
parameter signed W5TO34 = 0;
parameter signed W5TO35 = 0;
parameter signed W5TO36 = 0;
parameter signed W5TO37 = 0;
parameter signed W5TO38 = 0;
parameter signed W5TO39 = 0;
parameter signed W5TO40 = 0;
parameter signed W5TO41 = 0;
parameter signed W5TO42 = 0;
parameter signed W5TO43 = 0;
parameter signed W5TO44 = 0;
parameter signed W5TO45 = 0;
parameter signed W5TO46 = 0;
parameter signed W5TO47 = 0;
parameter signed W5TO48 = 0;
parameter signed W5TO49 = 0;
parameter signed W5TO50 = 0;
parameter signed W5TO51 = 0;
parameter signed W5TO52 = 0;
parameter signed W5TO53 = 0;
parameter signed W5TO54 = 0;
parameter signed W5TO55 = 0;
parameter signed W5TO56 = 0;
parameter signed W5TO57 = 0;
parameter signed W5TO58 = 0;
parameter signed W5TO59 = 0;
parameter signed W5TO60 = 0;
parameter signed W5TO61 = 0;
parameter signed W5TO62 = 0;
parameter signed W5TO63 = 0;
parameter signed W6TO0 = 0;
parameter signed W6TO1 = 0;
parameter signed W6TO2 = 0;
parameter signed W6TO3 = 0;
parameter signed W6TO4 = 0;
parameter signed W6TO5 = 0;
parameter signed W6TO6 = 0;
parameter signed W6TO7 = 0;
parameter signed W6TO8 = 0;
parameter signed W6TO9 = 0;
parameter signed W6TO10 = 0;
parameter signed W6TO11 = 0;
parameter signed W6TO12 = 0;
parameter signed W6TO13 = 0;
parameter signed W6TO14 = 0;
parameter signed W6TO15 = 0;
parameter signed W6TO16 = 0;
parameter signed W6TO17 = 0;
parameter signed W6TO18 = 0;
parameter signed W6TO19 = 0;
parameter signed W6TO20 = 0;
parameter signed W6TO21 = 0;
parameter signed W6TO22 = 0;
parameter signed W6TO23 = 0;
parameter signed W6TO24 = 0;
parameter signed W6TO25 = 0;
parameter signed W6TO26 = 0;
parameter signed W6TO27 = 0;
parameter signed W6TO28 = 0;
parameter signed W6TO29 = 0;
parameter signed W6TO30 = 0;
parameter signed W6TO31 = 0;
parameter signed W6TO32 = 0;
parameter signed W6TO33 = 0;
parameter signed W6TO34 = 0;
parameter signed W6TO35 = 0;
parameter signed W6TO36 = 0;
parameter signed W6TO37 = 0;
parameter signed W6TO38 = 0;
parameter signed W6TO39 = 0;
parameter signed W6TO40 = 0;
parameter signed W6TO41 = 0;
parameter signed W6TO42 = 0;
parameter signed W6TO43 = 0;
parameter signed W6TO44 = 0;
parameter signed W6TO45 = 0;
parameter signed W6TO46 = 0;
parameter signed W6TO47 = 0;
parameter signed W6TO48 = 0;
parameter signed W6TO49 = 0;
parameter signed W6TO50 = 0;
parameter signed W6TO51 = 0;
parameter signed W6TO52 = 0;
parameter signed W6TO53 = 0;
parameter signed W6TO54 = 0;
parameter signed W6TO55 = 0;
parameter signed W6TO56 = 0;
parameter signed W6TO57 = 0;
parameter signed W6TO58 = 0;
parameter signed W6TO59 = 0;
parameter signed W6TO60 = 0;
parameter signed W6TO61 = 0;
parameter signed W6TO62 = 0;
parameter signed W6TO63 = 0;
parameter signed W7TO0 = 0;
parameter signed W7TO1 = 0;
parameter signed W7TO2 = 0;
parameter signed W7TO3 = 0;
parameter signed W7TO4 = 0;
parameter signed W7TO5 = 0;
parameter signed W7TO6 = 0;
parameter signed W7TO7 = 0;
parameter signed W7TO8 = 0;
parameter signed W7TO9 = 0;
parameter signed W7TO10 = 0;
parameter signed W7TO11 = 0;
parameter signed W7TO12 = 0;
parameter signed W7TO13 = 0;
parameter signed W7TO14 = 0;
parameter signed W7TO15 = 0;
parameter signed W7TO16 = 0;
parameter signed W7TO17 = 0;
parameter signed W7TO18 = 0;
parameter signed W7TO19 = 0;
parameter signed W7TO20 = 0;
parameter signed W7TO21 = 0;
parameter signed W7TO22 = 0;
parameter signed W7TO23 = 0;
parameter signed W7TO24 = 0;
parameter signed W7TO25 = 0;
parameter signed W7TO26 = 0;
parameter signed W7TO27 = 0;
parameter signed W7TO28 = 0;
parameter signed W7TO29 = 0;
parameter signed W7TO30 = 0;
parameter signed W7TO31 = 0;
parameter signed W7TO32 = 0;
parameter signed W7TO33 = 0;
parameter signed W7TO34 = 0;
parameter signed W7TO35 = 0;
parameter signed W7TO36 = 0;
parameter signed W7TO37 = 0;
parameter signed W7TO38 = 0;
parameter signed W7TO39 = 0;
parameter signed W7TO40 = 0;
parameter signed W7TO41 = 0;
parameter signed W7TO42 = 0;
parameter signed W7TO43 = 0;
parameter signed W7TO44 = 0;
parameter signed W7TO45 = 0;
parameter signed W7TO46 = 0;
parameter signed W7TO47 = 0;
parameter signed W7TO48 = 0;
parameter signed W7TO49 = 0;
parameter signed W7TO50 = 0;
parameter signed W7TO51 = 0;
parameter signed W7TO52 = 0;
parameter signed W7TO53 = 0;
parameter signed W7TO54 = 0;
parameter signed W7TO55 = 0;
parameter signed W7TO56 = 0;
parameter signed W7TO57 = 0;
parameter signed W7TO58 = 0;
parameter signed W7TO59 = 0;
parameter signed W7TO60 = 0;
parameter signed W7TO61 = 0;
parameter signed W7TO62 = 0;
parameter signed W7TO63 = 0;
parameter signed W8TO0 = 0;
parameter signed W8TO1 = 0;
parameter signed W8TO2 = 0;
parameter signed W8TO3 = 0;
parameter signed W8TO4 = 0;
parameter signed W8TO5 = 0;
parameter signed W8TO6 = 0;
parameter signed W8TO7 = 0;
parameter signed W8TO8 = 0;
parameter signed W8TO9 = 0;
parameter signed W8TO10 = 0;
parameter signed W8TO11 = 0;
parameter signed W8TO12 = 0;
parameter signed W8TO13 = 0;
parameter signed W8TO14 = 0;
parameter signed W8TO15 = 0;
parameter signed W8TO16 = 0;
parameter signed W8TO17 = 0;
parameter signed W8TO18 = 0;
parameter signed W8TO19 = 0;
parameter signed W8TO20 = 0;
parameter signed W8TO21 = 0;
parameter signed W8TO22 = 0;
parameter signed W8TO23 = 0;
parameter signed W8TO24 = 0;
parameter signed W8TO25 = 0;
parameter signed W8TO26 = 0;
parameter signed W8TO27 = 0;
parameter signed W8TO28 = 0;
parameter signed W8TO29 = 0;
parameter signed W8TO30 = 0;
parameter signed W8TO31 = 0;
parameter signed W8TO32 = 0;
parameter signed W8TO33 = 0;
parameter signed W8TO34 = 0;
parameter signed W8TO35 = 0;
parameter signed W8TO36 = 0;
parameter signed W8TO37 = 0;
parameter signed W8TO38 = 0;
parameter signed W8TO39 = 0;
parameter signed W8TO40 = 0;
parameter signed W8TO41 = 0;
parameter signed W8TO42 = 0;
parameter signed W8TO43 = 0;
parameter signed W8TO44 = 0;
parameter signed W8TO45 = 0;
parameter signed W8TO46 = 0;
parameter signed W8TO47 = 0;
parameter signed W8TO48 = 0;
parameter signed W8TO49 = 0;
parameter signed W8TO50 = 0;
parameter signed W8TO51 = 0;
parameter signed W8TO52 = 0;
parameter signed W8TO53 = 0;
parameter signed W8TO54 = 0;
parameter signed W8TO55 = 0;
parameter signed W8TO56 = 0;
parameter signed W8TO57 = 0;
parameter signed W8TO58 = 0;
parameter signed W8TO59 = 0;
parameter signed W8TO60 = 0;
parameter signed W8TO61 = 0;
parameter signed W8TO62 = 0;
parameter signed W8TO63 = 0;
parameter signed W9TO0 = 0;
parameter signed W9TO1 = 0;
parameter signed W9TO2 = 0;
parameter signed W9TO3 = 0;
parameter signed W9TO4 = 0;
parameter signed W9TO5 = 0;
parameter signed W9TO6 = 0;
parameter signed W9TO7 = 0;
parameter signed W9TO8 = 0;
parameter signed W9TO9 = 0;
parameter signed W9TO10 = 0;
parameter signed W9TO11 = 0;
parameter signed W9TO12 = 0;
parameter signed W9TO13 = 0;
parameter signed W9TO14 = 0;
parameter signed W9TO15 = 0;
parameter signed W9TO16 = 0;
parameter signed W9TO17 = 0;
parameter signed W9TO18 = 0;
parameter signed W9TO19 = 0;
parameter signed W9TO20 = 0;
parameter signed W9TO21 = 0;
parameter signed W9TO22 = 0;
parameter signed W9TO23 = 0;
parameter signed W9TO24 = 0;
parameter signed W9TO25 = 0;
parameter signed W9TO26 = 0;
parameter signed W9TO27 = 0;
parameter signed W9TO28 = 0;
parameter signed W9TO29 = 0;
parameter signed W9TO30 = 0;
parameter signed W9TO31 = 0;
parameter signed W9TO32 = 0;
parameter signed W9TO33 = 0;
parameter signed W9TO34 = 0;
parameter signed W9TO35 = 0;
parameter signed W9TO36 = 0;
parameter signed W9TO37 = 0;
parameter signed W9TO38 = 0;
parameter signed W9TO39 = 0;
parameter signed W9TO40 = 0;
parameter signed W9TO41 = 0;
parameter signed W9TO42 = 0;
parameter signed W9TO43 = 0;
parameter signed W9TO44 = 0;
parameter signed W9TO45 = 0;
parameter signed W9TO46 = 0;
parameter signed W9TO47 = 0;
parameter signed W9TO48 = 0;
parameter signed W9TO49 = 0;
parameter signed W9TO50 = 0;
parameter signed W9TO51 = 0;
parameter signed W9TO52 = 0;
parameter signed W9TO53 = 0;
parameter signed W9TO54 = 0;
parameter signed W9TO55 = 0;
parameter signed W9TO56 = 0;
parameter signed W9TO57 = 0;
parameter signed W9TO58 = 0;
parameter signed W9TO59 = 0;
parameter signed W9TO60 = 0;
parameter signed W9TO61 = 0;
parameter signed W9TO62 = 0;
parameter signed W9TO63 = 0;
parameter signed W10TO0 = 0;
parameter signed W10TO1 = 0;
parameter signed W10TO2 = 0;
parameter signed W10TO3 = 0;
parameter signed W10TO4 = 0;
parameter signed W10TO5 = 0;
parameter signed W10TO6 = 0;
parameter signed W10TO7 = 0;
parameter signed W10TO8 = 0;
parameter signed W10TO9 = 0;
parameter signed W10TO10 = 0;
parameter signed W10TO11 = 0;
parameter signed W10TO12 = 0;
parameter signed W10TO13 = 0;
parameter signed W10TO14 = 0;
parameter signed W10TO15 = 0;
parameter signed W10TO16 = 0;
parameter signed W10TO17 = 0;
parameter signed W10TO18 = 0;
parameter signed W10TO19 = 0;
parameter signed W10TO20 = 0;
parameter signed W10TO21 = 0;
parameter signed W10TO22 = 0;
parameter signed W10TO23 = 0;
parameter signed W10TO24 = 0;
parameter signed W10TO25 = 0;
parameter signed W10TO26 = 0;
parameter signed W10TO27 = 0;
parameter signed W10TO28 = 0;
parameter signed W10TO29 = 0;
parameter signed W10TO30 = 0;
parameter signed W10TO31 = 0;
parameter signed W10TO32 = 0;
parameter signed W10TO33 = 0;
parameter signed W10TO34 = 0;
parameter signed W10TO35 = 0;
parameter signed W10TO36 = 0;
parameter signed W10TO37 = 0;
parameter signed W10TO38 = 0;
parameter signed W10TO39 = 0;
parameter signed W10TO40 = 0;
parameter signed W10TO41 = 0;
parameter signed W10TO42 = 0;
parameter signed W10TO43 = 0;
parameter signed W10TO44 = 0;
parameter signed W10TO45 = 0;
parameter signed W10TO46 = 0;
parameter signed W10TO47 = 0;
parameter signed W10TO48 = 0;
parameter signed W10TO49 = 0;
parameter signed W10TO50 = 0;
parameter signed W10TO51 = 0;
parameter signed W10TO52 = 0;
parameter signed W10TO53 = 0;
parameter signed W10TO54 = 0;
parameter signed W10TO55 = 0;
parameter signed W10TO56 = 0;
parameter signed W10TO57 = 0;
parameter signed W10TO58 = 0;
parameter signed W10TO59 = 0;
parameter signed W10TO60 = 0;
parameter signed W10TO61 = 0;
parameter signed W10TO62 = 0;
parameter signed W10TO63 = 0;
parameter signed W11TO0 = 0;
parameter signed W11TO1 = 0;
parameter signed W11TO2 = 0;
parameter signed W11TO3 = 0;
parameter signed W11TO4 = 0;
parameter signed W11TO5 = 0;
parameter signed W11TO6 = 0;
parameter signed W11TO7 = 0;
parameter signed W11TO8 = 0;
parameter signed W11TO9 = 0;
parameter signed W11TO10 = 0;
parameter signed W11TO11 = 0;
parameter signed W11TO12 = 0;
parameter signed W11TO13 = 0;
parameter signed W11TO14 = 0;
parameter signed W11TO15 = 0;
parameter signed W11TO16 = 0;
parameter signed W11TO17 = 0;
parameter signed W11TO18 = 0;
parameter signed W11TO19 = 0;
parameter signed W11TO20 = 0;
parameter signed W11TO21 = 0;
parameter signed W11TO22 = 0;
parameter signed W11TO23 = 0;
parameter signed W11TO24 = 0;
parameter signed W11TO25 = 0;
parameter signed W11TO26 = 0;
parameter signed W11TO27 = 0;
parameter signed W11TO28 = 0;
parameter signed W11TO29 = 0;
parameter signed W11TO30 = 0;
parameter signed W11TO31 = 0;
parameter signed W11TO32 = 0;
parameter signed W11TO33 = 0;
parameter signed W11TO34 = 0;
parameter signed W11TO35 = 0;
parameter signed W11TO36 = 0;
parameter signed W11TO37 = 0;
parameter signed W11TO38 = 0;
parameter signed W11TO39 = 0;
parameter signed W11TO40 = 0;
parameter signed W11TO41 = 0;
parameter signed W11TO42 = 0;
parameter signed W11TO43 = 0;
parameter signed W11TO44 = 0;
parameter signed W11TO45 = 0;
parameter signed W11TO46 = 0;
parameter signed W11TO47 = 0;
parameter signed W11TO48 = 0;
parameter signed W11TO49 = 0;
parameter signed W11TO50 = 0;
parameter signed W11TO51 = 0;
parameter signed W11TO52 = 0;
parameter signed W11TO53 = 0;
parameter signed W11TO54 = 0;
parameter signed W11TO55 = 0;
parameter signed W11TO56 = 0;
parameter signed W11TO57 = 0;
parameter signed W11TO58 = 0;
parameter signed W11TO59 = 0;
parameter signed W11TO60 = 0;
parameter signed W11TO61 = 0;
parameter signed W11TO62 = 0;
parameter signed W11TO63 = 0;
parameter signed W12TO0 = 0;
parameter signed W12TO1 = 0;
parameter signed W12TO2 = 0;
parameter signed W12TO3 = 0;
parameter signed W12TO4 = 0;
parameter signed W12TO5 = 0;
parameter signed W12TO6 = 0;
parameter signed W12TO7 = 0;
parameter signed W12TO8 = 0;
parameter signed W12TO9 = 0;
parameter signed W12TO10 = 0;
parameter signed W12TO11 = 0;
parameter signed W12TO12 = 0;
parameter signed W12TO13 = 0;
parameter signed W12TO14 = 0;
parameter signed W12TO15 = 0;
parameter signed W12TO16 = 0;
parameter signed W12TO17 = 0;
parameter signed W12TO18 = 0;
parameter signed W12TO19 = 0;
parameter signed W12TO20 = 0;
parameter signed W12TO21 = 0;
parameter signed W12TO22 = 0;
parameter signed W12TO23 = 0;
parameter signed W12TO24 = 0;
parameter signed W12TO25 = 0;
parameter signed W12TO26 = 0;
parameter signed W12TO27 = 0;
parameter signed W12TO28 = 0;
parameter signed W12TO29 = 0;
parameter signed W12TO30 = 0;
parameter signed W12TO31 = 0;
parameter signed W12TO32 = 0;
parameter signed W12TO33 = 0;
parameter signed W12TO34 = 0;
parameter signed W12TO35 = 0;
parameter signed W12TO36 = 0;
parameter signed W12TO37 = 0;
parameter signed W12TO38 = 0;
parameter signed W12TO39 = 0;
parameter signed W12TO40 = 0;
parameter signed W12TO41 = 0;
parameter signed W12TO42 = 0;
parameter signed W12TO43 = 0;
parameter signed W12TO44 = 0;
parameter signed W12TO45 = 0;
parameter signed W12TO46 = 0;
parameter signed W12TO47 = 0;
parameter signed W12TO48 = 0;
parameter signed W12TO49 = 0;
parameter signed W12TO50 = 0;
parameter signed W12TO51 = 0;
parameter signed W12TO52 = 0;
parameter signed W12TO53 = 0;
parameter signed W12TO54 = 0;
parameter signed W12TO55 = 0;
parameter signed W12TO56 = 0;
parameter signed W12TO57 = 0;
parameter signed W12TO58 = 0;
parameter signed W12TO59 = 0;
parameter signed W12TO60 = 0;
parameter signed W12TO61 = 0;
parameter signed W12TO62 = 0;
parameter signed W12TO63 = 0;
parameter signed W13TO0 = 0;
parameter signed W13TO1 = 0;
parameter signed W13TO2 = 0;
parameter signed W13TO3 = 0;
parameter signed W13TO4 = 0;
parameter signed W13TO5 = 0;
parameter signed W13TO6 = 0;
parameter signed W13TO7 = 0;
parameter signed W13TO8 = 0;
parameter signed W13TO9 = 0;
parameter signed W13TO10 = 0;
parameter signed W13TO11 = 0;
parameter signed W13TO12 = 0;
parameter signed W13TO13 = 0;
parameter signed W13TO14 = 0;
parameter signed W13TO15 = 0;
parameter signed W13TO16 = 0;
parameter signed W13TO17 = 0;
parameter signed W13TO18 = 0;
parameter signed W13TO19 = 0;
parameter signed W13TO20 = 0;
parameter signed W13TO21 = 0;
parameter signed W13TO22 = 0;
parameter signed W13TO23 = 0;
parameter signed W13TO24 = 0;
parameter signed W13TO25 = 0;
parameter signed W13TO26 = 0;
parameter signed W13TO27 = 0;
parameter signed W13TO28 = 0;
parameter signed W13TO29 = 0;
parameter signed W13TO30 = 0;
parameter signed W13TO31 = 0;
parameter signed W13TO32 = 0;
parameter signed W13TO33 = 0;
parameter signed W13TO34 = 0;
parameter signed W13TO35 = 0;
parameter signed W13TO36 = 0;
parameter signed W13TO37 = 0;
parameter signed W13TO38 = 0;
parameter signed W13TO39 = 0;
parameter signed W13TO40 = 0;
parameter signed W13TO41 = 0;
parameter signed W13TO42 = 0;
parameter signed W13TO43 = 0;
parameter signed W13TO44 = 0;
parameter signed W13TO45 = 0;
parameter signed W13TO46 = 0;
parameter signed W13TO47 = 0;
parameter signed W13TO48 = 0;
parameter signed W13TO49 = 0;
parameter signed W13TO50 = 0;
parameter signed W13TO51 = 0;
parameter signed W13TO52 = 0;
parameter signed W13TO53 = 0;
parameter signed W13TO54 = 0;
parameter signed W13TO55 = 0;
parameter signed W13TO56 = 0;
parameter signed W13TO57 = 0;
parameter signed W13TO58 = 0;
parameter signed W13TO59 = 0;
parameter signed W13TO60 = 0;
parameter signed W13TO61 = 0;
parameter signed W13TO62 = 0;
parameter signed W13TO63 = 0;
parameter signed W14TO0 = 0;
parameter signed W14TO1 = 0;
parameter signed W14TO2 = 0;
parameter signed W14TO3 = 0;
parameter signed W14TO4 = 0;
parameter signed W14TO5 = 0;
parameter signed W14TO6 = 0;
parameter signed W14TO7 = 0;
parameter signed W14TO8 = 0;
parameter signed W14TO9 = 0;
parameter signed W14TO10 = 0;
parameter signed W14TO11 = 0;
parameter signed W14TO12 = 0;
parameter signed W14TO13 = 0;
parameter signed W14TO14 = 0;
parameter signed W14TO15 = 0;
parameter signed W14TO16 = 0;
parameter signed W14TO17 = 0;
parameter signed W14TO18 = 0;
parameter signed W14TO19 = 0;
parameter signed W14TO20 = 0;
parameter signed W14TO21 = 0;
parameter signed W14TO22 = 0;
parameter signed W14TO23 = 0;
parameter signed W14TO24 = 0;
parameter signed W14TO25 = 0;
parameter signed W14TO26 = 0;
parameter signed W14TO27 = 0;
parameter signed W14TO28 = 0;
parameter signed W14TO29 = 0;
parameter signed W14TO30 = 0;
parameter signed W14TO31 = 0;
parameter signed W14TO32 = 0;
parameter signed W14TO33 = 0;
parameter signed W14TO34 = 0;
parameter signed W14TO35 = 0;
parameter signed W14TO36 = 0;
parameter signed W14TO37 = 0;
parameter signed W14TO38 = 0;
parameter signed W14TO39 = 0;
parameter signed W14TO40 = 0;
parameter signed W14TO41 = 0;
parameter signed W14TO42 = 0;
parameter signed W14TO43 = 0;
parameter signed W14TO44 = 0;
parameter signed W14TO45 = 0;
parameter signed W14TO46 = 0;
parameter signed W14TO47 = 0;
parameter signed W14TO48 = 0;
parameter signed W14TO49 = 0;
parameter signed W14TO50 = 0;
parameter signed W14TO51 = 0;
parameter signed W14TO52 = 0;
parameter signed W14TO53 = 0;
parameter signed W14TO54 = 0;
parameter signed W14TO55 = 0;
parameter signed W14TO56 = 0;
parameter signed W14TO57 = 0;
parameter signed W14TO58 = 0;
parameter signed W14TO59 = 0;
parameter signed W14TO60 = 0;
parameter signed W14TO61 = 0;
parameter signed W14TO62 = 0;
parameter signed W14TO63 = 0;
parameter signed W15TO0 = 0;
parameter signed W15TO1 = 0;
parameter signed W15TO2 = 0;
parameter signed W15TO3 = 0;
parameter signed W15TO4 = 0;
parameter signed W15TO5 = 0;
parameter signed W15TO6 = 0;
parameter signed W15TO7 = 0;
parameter signed W15TO8 = 0;
parameter signed W15TO9 = 0;
parameter signed W15TO10 = 0;
parameter signed W15TO11 = 0;
parameter signed W15TO12 = 0;
parameter signed W15TO13 = 0;
parameter signed W15TO14 = 0;
parameter signed W15TO15 = 0;
parameter signed W15TO16 = 0;
parameter signed W15TO17 = 0;
parameter signed W15TO18 = 0;
parameter signed W15TO19 = 0;
parameter signed W15TO20 = 0;
parameter signed W15TO21 = 0;
parameter signed W15TO22 = 0;
parameter signed W15TO23 = 0;
parameter signed W15TO24 = 0;
parameter signed W15TO25 = 0;
parameter signed W15TO26 = 0;
parameter signed W15TO27 = 0;
parameter signed W15TO28 = 0;
parameter signed W15TO29 = 0;
parameter signed W15TO30 = 0;
parameter signed W15TO31 = 0;
parameter signed W15TO32 = 0;
parameter signed W15TO33 = 0;
parameter signed W15TO34 = 0;
parameter signed W15TO35 = 0;
parameter signed W15TO36 = 0;
parameter signed W15TO37 = 0;
parameter signed W15TO38 = 0;
parameter signed W15TO39 = 0;
parameter signed W15TO40 = 0;
parameter signed W15TO41 = 0;
parameter signed W15TO42 = 0;
parameter signed W15TO43 = 0;
parameter signed W15TO44 = 0;
parameter signed W15TO45 = 0;
parameter signed W15TO46 = 0;
parameter signed W15TO47 = 0;
parameter signed W15TO48 = 0;
parameter signed W15TO49 = 0;
parameter signed W15TO50 = 0;
parameter signed W15TO51 = 0;
parameter signed W15TO52 = 0;
parameter signed W15TO53 = 0;
parameter signed W15TO54 = 0;
parameter signed W15TO55 = 0;
parameter signed W15TO56 = 0;
parameter signed W15TO57 = 0;
parameter signed W15TO58 = 0;
parameter signed W15TO59 = 0;
parameter signed W15TO60 = 0;
parameter signed W15TO61 = 0;
parameter signed W15TO62 = 0;
parameter signed W15TO63 = 0;
parameter signed W16TO0 = 0;
parameter signed W16TO1 = 0;
parameter signed W16TO2 = 0;
parameter signed W16TO3 = 0;
parameter signed W16TO4 = 0;
parameter signed W16TO5 = 0;
parameter signed W16TO6 = 0;
parameter signed W16TO7 = 0;
parameter signed W16TO8 = 0;
parameter signed W16TO9 = 0;
parameter signed W16TO10 = 0;
parameter signed W16TO11 = 0;
parameter signed W16TO12 = 0;
parameter signed W16TO13 = 0;
parameter signed W16TO14 = 0;
parameter signed W16TO15 = 0;
parameter signed W16TO16 = 0;
parameter signed W16TO17 = 0;
parameter signed W16TO18 = 0;
parameter signed W16TO19 = 0;
parameter signed W16TO20 = 0;
parameter signed W16TO21 = 0;
parameter signed W16TO22 = 0;
parameter signed W16TO23 = 0;
parameter signed W16TO24 = 0;
parameter signed W16TO25 = 0;
parameter signed W16TO26 = 0;
parameter signed W16TO27 = 0;
parameter signed W16TO28 = 0;
parameter signed W16TO29 = 0;
parameter signed W16TO30 = 0;
parameter signed W16TO31 = 0;
parameter signed W16TO32 = 0;
parameter signed W16TO33 = 0;
parameter signed W16TO34 = 0;
parameter signed W16TO35 = 0;
parameter signed W16TO36 = 0;
parameter signed W16TO37 = 0;
parameter signed W16TO38 = 0;
parameter signed W16TO39 = 0;
parameter signed W16TO40 = 0;
parameter signed W16TO41 = 0;
parameter signed W16TO42 = 0;
parameter signed W16TO43 = 0;
parameter signed W16TO44 = 0;
parameter signed W16TO45 = 0;
parameter signed W16TO46 = 0;
parameter signed W16TO47 = 0;
parameter signed W16TO48 = 0;
parameter signed W16TO49 = 0;
parameter signed W16TO50 = 0;
parameter signed W16TO51 = 0;
parameter signed W16TO52 = 0;
parameter signed W16TO53 = 0;
parameter signed W16TO54 = 0;
parameter signed W16TO55 = 0;
parameter signed W16TO56 = 0;
parameter signed W16TO57 = 0;
parameter signed W16TO58 = 0;
parameter signed W16TO59 = 0;
parameter signed W16TO60 = 0;
parameter signed W16TO61 = 0;
parameter signed W16TO62 = 0;
parameter signed W16TO63 = 0;
parameter signed W17TO0 = 0;
parameter signed W17TO1 = 0;
parameter signed W17TO2 = 0;
parameter signed W17TO3 = 0;
parameter signed W17TO4 = 0;
parameter signed W17TO5 = 0;
parameter signed W17TO6 = 0;
parameter signed W17TO7 = 0;
parameter signed W17TO8 = 0;
parameter signed W17TO9 = 0;
parameter signed W17TO10 = 0;
parameter signed W17TO11 = 0;
parameter signed W17TO12 = 0;
parameter signed W17TO13 = 0;
parameter signed W17TO14 = 0;
parameter signed W17TO15 = 0;
parameter signed W17TO16 = 0;
parameter signed W17TO17 = 0;
parameter signed W17TO18 = 0;
parameter signed W17TO19 = 0;
parameter signed W17TO20 = 0;
parameter signed W17TO21 = 0;
parameter signed W17TO22 = 0;
parameter signed W17TO23 = 0;
parameter signed W17TO24 = 0;
parameter signed W17TO25 = 0;
parameter signed W17TO26 = 0;
parameter signed W17TO27 = 0;
parameter signed W17TO28 = 0;
parameter signed W17TO29 = 0;
parameter signed W17TO30 = 0;
parameter signed W17TO31 = 0;
parameter signed W17TO32 = 0;
parameter signed W17TO33 = 0;
parameter signed W17TO34 = 0;
parameter signed W17TO35 = 0;
parameter signed W17TO36 = 0;
parameter signed W17TO37 = 0;
parameter signed W17TO38 = 0;
parameter signed W17TO39 = 0;
parameter signed W17TO40 = 0;
parameter signed W17TO41 = 0;
parameter signed W17TO42 = 0;
parameter signed W17TO43 = 0;
parameter signed W17TO44 = 0;
parameter signed W17TO45 = 0;
parameter signed W17TO46 = 0;
parameter signed W17TO47 = 0;
parameter signed W17TO48 = 0;
parameter signed W17TO49 = 0;
parameter signed W17TO50 = 0;
parameter signed W17TO51 = 0;
parameter signed W17TO52 = 0;
parameter signed W17TO53 = 0;
parameter signed W17TO54 = 0;
parameter signed W17TO55 = 0;
parameter signed W17TO56 = 0;
parameter signed W17TO57 = 0;
parameter signed W17TO58 = 0;
parameter signed W17TO59 = 0;
parameter signed W17TO60 = 0;
parameter signed W17TO61 = 0;
parameter signed W17TO62 = 0;
parameter signed W17TO63 = 0;
parameter signed W18TO0 = 0;
parameter signed W18TO1 = 0;
parameter signed W18TO2 = 0;
parameter signed W18TO3 = 0;
parameter signed W18TO4 = 0;
parameter signed W18TO5 = 0;
parameter signed W18TO6 = 0;
parameter signed W18TO7 = 0;
parameter signed W18TO8 = 0;
parameter signed W18TO9 = 0;
parameter signed W18TO10 = 0;
parameter signed W18TO11 = 0;
parameter signed W18TO12 = 0;
parameter signed W18TO13 = 0;
parameter signed W18TO14 = 0;
parameter signed W18TO15 = 0;
parameter signed W18TO16 = 0;
parameter signed W18TO17 = 0;
parameter signed W18TO18 = 0;
parameter signed W18TO19 = 0;
parameter signed W18TO20 = 0;
parameter signed W18TO21 = 0;
parameter signed W18TO22 = 0;
parameter signed W18TO23 = 0;
parameter signed W18TO24 = 0;
parameter signed W18TO25 = 0;
parameter signed W18TO26 = 0;
parameter signed W18TO27 = 0;
parameter signed W18TO28 = 0;
parameter signed W18TO29 = 0;
parameter signed W18TO30 = 0;
parameter signed W18TO31 = 0;
parameter signed W18TO32 = 0;
parameter signed W18TO33 = 0;
parameter signed W18TO34 = 0;
parameter signed W18TO35 = 0;
parameter signed W18TO36 = 0;
parameter signed W18TO37 = 0;
parameter signed W18TO38 = 0;
parameter signed W18TO39 = 0;
parameter signed W18TO40 = 0;
parameter signed W18TO41 = 0;
parameter signed W18TO42 = 0;
parameter signed W18TO43 = 0;
parameter signed W18TO44 = 0;
parameter signed W18TO45 = 0;
parameter signed W18TO46 = 0;
parameter signed W18TO47 = 0;
parameter signed W18TO48 = 0;
parameter signed W18TO49 = 0;
parameter signed W18TO50 = 0;
parameter signed W18TO51 = 0;
parameter signed W18TO52 = 0;
parameter signed W18TO53 = 0;
parameter signed W18TO54 = 0;
parameter signed W18TO55 = 0;
parameter signed W18TO56 = 0;
parameter signed W18TO57 = 0;
parameter signed W18TO58 = 0;
parameter signed W18TO59 = 0;
parameter signed W18TO60 = 0;
parameter signed W18TO61 = 0;
parameter signed W18TO62 = 0;
parameter signed W18TO63 = 0;
parameter signed W19TO0 = 0;
parameter signed W19TO1 = 0;
parameter signed W19TO2 = 0;
parameter signed W19TO3 = 0;
parameter signed W19TO4 = 0;
parameter signed W19TO5 = 0;
parameter signed W19TO6 = 0;
parameter signed W19TO7 = 0;
parameter signed W19TO8 = 0;
parameter signed W19TO9 = 0;
parameter signed W19TO10 = 0;
parameter signed W19TO11 = 0;
parameter signed W19TO12 = 0;
parameter signed W19TO13 = 0;
parameter signed W19TO14 = 0;
parameter signed W19TO15 = 0;
parameter signed W19TO16 = 0;
parameter signed W19TO17 = 0;
parameter signed W19TO18 = 0;
parameter signed W19TO19 = 0;
parameter signed W19TO20 = 0;
parameter signed W19TO21 = 0;
parameter signed W19TO22 = 0;
parameter signed W19TO23 = 0;
parameter signed W19TO24 = 0;
parameter signed W19TO25 = 0;
parameter signed W19TO26 = 0;
parameter signed W19TO27 = 0;
parameter signed W19TO28 = 0;
parameter signed W19TO29 = 0;
parameter signed W19TO30 = 0;
parameter signed W19TO31 = 0;
parameter signed W19TO32 = 0;
parameter signed W19TO33 = 0;
parameter signed W19TO34 = 0;
parameter signed W19TO35 = 0;
parameter signed W19TO36 = 0;
parameter signed W19TO37 = 0;
parameter signed W19TO38 = 0;
parameter signed W19TO39 = 0;
parameter signed W19TO40 = 0;
parameter signed W19TO41 = 0;
parameter signed W19TO42 = 0;
parameter signed W19TO43 = 0;
parameter signed W19TO44 = 0;
parameter signed W19TO45 = 0;
parameter signed W19TO46 = 0;
parameter signed W19TO47 = 0;
parameter signed W19TO48 = 0;
parameter signed W19TO49 = 0;
parameter signed W19TO50 = 0;
parameter signed W19TO51 = 0;
parameter signed W19TO52 = 0;
parameter signed W19TO53 = 0;
parameter signed W19TO54 = 0;
parameter signed W19TO55 = 0;
parameter signed W19TO56 = 0;
parameter signed W19TO57 = 0;
parameter signed W19TO58 = 0;
parameter signed W19TO59 = 0;
parameter signed W19TO60 = 0;
parameter signed W19TO61 = 0;
parameter signed W19TO62 = 0;
parameter signed W19TO63 = 0;
parameter signed W20TO0 = 0;
parameter signed W20TO1 = 0;
parameter signed W20TO2 = 0;
parameter signed W20TO3 = 0;
parameter signed W20TO4 = 0;
parameter signed W20TO5 = 0;
parameter signed W20TO6 = 0;
parameter signed W20TO7 = 0;
parameter signed W20TO8 = 0;
parameter signed W20TO9 = 0;
parameter signed W20TO10 = 0;
parameter signed W20TO11 = 0;
parameter signed W20TO12 = 0;
parameter signed W20TO13 = 0;
parameter signed W20TO14 = 0;
parameter signed W20TO15 = 0;
parameter signed W20TO16 = 0;
parameter signed W20TO17 = 0;
parameter signed W20TO18 = 0;
parameter signed W20TO19 = 0;
parameter signed W20TO20 = 0;
parameter signed W20TO21 = 0;
parameter signed W20TO22 = 0;
parameter signed W20TO23 = 0;
parameter signed W20TO24 = 0;
parameter signed W20TO25 = 0;
parameter signed W20TO26 = 0;
parameter signed W20TO27 = 0;
parameter signed W20TO28 = 0;
parameter signed W20TO29 = 0;
parameter signed W20TO30 = 0;
parameter signed W20TO31 = 0;
parameter signed W20TO32 = 0;
parameter signed W20TO33 = 0;
parameter signed W20TO34 = 0;
parameter signed W20TO35 = 0;
parameter signed W20TO36 = 0;
parameter signed W20TO37 = 0;
parameter signed W20TO38 = 0;
parameter signed W20TO39 = 0;
parameter signed W20TO40 = 0;
parameter signed W20TO41 = 0;
parameter signed W20TO42 = 0;
parameter signed W20TO43 = 0;
parameter signed W20TO44 = 0;
parameter signed W20TO45 = 0;
parameter signed W20TO46 = 0;
parameter signed W20TO47 = 0;
parameter signed W20TO48 = 0;
parameter signed W20TO49 = 0;
parameter signed W20TO50 = 0;
parameter signed W20TO51 = 0;
parameter signed W20TO52 = 0;
parameter signed W20TO53 = 0;
parameter signed W20TO54 = 0;
parameter signed W20TO55 = 0;
parameter signed W20TO56 = 0;
parameter signed W20TO57 = 0;
parameter signed W20TO58 = 0;
parameter signed W20TO59 = 0;
parameter signed W20TO60 = 0;
parameter signed W20TO61 = 0;
parameter signed W20TO62 = 0;
parameter signed W20TO63 = 0;
parameter signed W21TO0 = 0;
parameter signed W21TO1 = 0;
parameter signed W21TO2 = 0;
parameter signed W21TO3 = 0;
parameter signed W21TO4 = 0;
parameter signed W21TO5 = 0;
parameter signed W21TO6 = 0;
parameter signed W21TO7 = 0;
parameter signed W21TO8 = 0;
parameter signed W21TO9 = 0;
parameter signed W21TO10 = 0;
parameter signed W21TO11 = 0;
parameter signed W21TO12 = 0;
parameter signed W21TO13 = 0;
parameter signed W21TO14 = 0;
parameter signed W21TO15 = 0;
parameter signed W21TO16 = 0;
parameter signed W21TO17 = 0;
parameter signed W21TO18 = 0;
parameter signed W21TO19 = 0;
parameter signed W21TO20 = 0;
parameter signed W21TO21 = 0;
parameter signed W21TO22 = 0;
parameter signed W21TO23 = 0;
parameter signed W21TO24 = 0;
parameter signed W21TO25 = 0;
parameter signed W21TO26 = 0;
parameter signed W21TO27 = 0;
parameter signed W21TO28 = 0;
parameter signed W21TO29 = 0;
parameter signed W21TO30 = 0;
parameter signed W21TO31 = 0;
parameter signed W21TO32 = 0;
parameter signed W21TO33 = 0;
parameter signed W21TO34 = 0;
parameter signed W21TO35 = 0;
parameter signed W21TO36 = 0;
parameter signed W21TO37 = 0;
parameter signed W21TO38 = 0;
parameter signed W21TO39 = 0;
parameter signed W21TO40 = 0;
parameter signed W21TO41 = 0;
parameter signed W21TO42 = 0;
parameter signed W21TO43 = 0;
parameter signed W21TO44 = 0;
parameter signed W21TO45 = 0;
parameter signed W21TO46 = 0;
parameter signed W21TO47 = 0;
parameter signed W21TO48 = 0;
parameter signed W21TO49 = 0;
parameter signed W21TO50 = 0;
parameter signed W21TO51 = 0;
parameter signed W21TO52 = 0;
parameter signed W21TO53 = 0;
parameter signed W21TO54 = 0;
parameter signed W21TO55 = 0;
parameter signed W21TO56 = 0;
parameter signed W21TO57 = 0;
parameter signed W21TO58 = 0;
parameter signed W21TO59 = 0;
parameter signed W21TO60 = 0;
parameter signed W21TO61 = 0;
parameter signed W21TO62 = 0;
parameter signed W21TO63 = 0;
parameter signed W22TO0 = 0;
parameter signed W22TO1 = 0;
parameter signed W22TO2 = 0;
parameter signed W22TO3 = 0;
parameter signed W22TO4 = 0;
parameter signed W22TO5 = 0;
parameter signed W22TO6 = 0;
parameter signed W22TO7 = 0;
parameter signed W22TO8 = 0;
parameter signed W22TO9 = 0;
parameter signed W22TO10 = 0;
parameter signed W22TO11 = 0;
parameter signed W22TO12 = 0;
parameter signed W22TO13 = 0;
parameter signed W22TO14 = 0;
parameter signed W22TO15 = 0;
parameter signed W22TO16 = 0;
parameter signed W22TO17 = 0;
parameter signed W22TO18 = 0;
parameter signed W22TO19 = 0;
parameter signed W22TO20 = 0;
parameter signed W22TO21 = 0;
parameter signed W22TO22 = 0;
parameter signed W22TO23 = 0;
parameter signed W22TO24 = 0;
parameter signed W22TO25 = 0;
parameter signed W22TO26 = 0;
parameter signed W22TO27 = 0;
parameter signed W22TO28 = 0;
parameter signed W22TO29 = 0;
parameter signed W22TO30 = 0;
parameter signed W22TO31 = 0;
parameter signed W22TO32 = 0;
parameter signed W22TO33 = 0;
parameter signed W22TO34 = 0;
parameter signed W22TO35 = 0;
parameter signed W22TO36 = 0;
parameter signed W22TO37 = 0;
parameter signed W22TO38 = 0;
parameter signed W22TO39 = 0;
parameter signed W22TO40 = 0;
parameter signed W22TO41 = 0;
parameter signed W22TO42 = 0;
parameter signed W22TO43 = 0;
parameter signed W22TO44 = 0;
parameter signed W22TO45 = 0;
parameter signed W22TO46 = 0;
parameter signed W22TO47 = 0;
parameter signed W22TO48 = 0;
parameter signed W22TO49 = 0;
parameter signed W22TO50 = 0;
parameter signed W22TO51 = 0;
parameter signed W22TO52 = 0;
parameter signed W22TO53 = 0;
parameter signed W22TO54 = 0;
parameter signed W22TO55 = 0;
parameter signed W22TO56 = 0;
parameter signed W22TO57 = 0;
parameter signed W22TO58 = 0;
parameter signed W22TO59 = 0;
parameter signed W22TO60 = 0;
parameter signed W22TO61 = 0;
parameter signed W22TO62 = 0;
parameter signed W22TO63 = 0;
parameter signed W23TO0 = 0;
parameter signed W23TO1 = 0;
parameter signed W23TO2 = 0;
parameter signed W23TO3 = 0;
parameter signed W23TO4 = 0;
parameter signed W23TO5 = 0;
parameter signed W23TO6 = 0;
parameter signed W23TO7 = 0;
parameter signed W23TO8 = 0;
parameter signed W23TO9 = 0;
parameter signed W23TO10 = 0;
parameter signed W23TO11 = 0;
parameter signed W23TO12 = 0;
parameter signed W23TO13 = 0;
parameter signed W23TO14 = 0;
parameter signed W23TO15 = 0;
parameter signed W23TO16 = 0;
parameter signed W23TO17 = 0;
parameter signed W23TO18 = 0;
parameter signed W23TO19 = 0;
parameter signed W23TO20 = 0;
parameter signed W23TO21 = 0;
parameter signed W23TO22 = 0;
parameter signed W23TO23 = 0;
parameter signed W23TO24 = 0;
parameter signed W23TO25 = 0;
parameter signed W23TO26 = 0;
parameter signed W23TO27 = 0;
parameter signed W23TO28 = 0;
parameter signed W23TO29 = 0;
parameter signed W23TO30 = 0;
parameter signed W23TO31 = 0;
parameter signed W23TO32 = 0;
parameter signed W23TO33 = 0;
parameter signed W23TO34 = 0;
parameter signed W23TO35 = 0;
parameter signed W23TO36 = 0;
parameter signed W23TO37 = 0;
parameter signed W23TO38 = 0;
parameter signed W23TO39 = 0;
parameter signed W23TO40 = 0;
parameter signed W23TO41 = 0;
parameter signed W23TO42 = 0;
parameter signed W23TO43 = 0;
parameter signed W23TO44 = 0;
parameter signed W23TO45 = 0;
parameter signed W23TO46 = 0;
parameter signed W23TO47 = 0;
parameter signed W23TO48 = 0;
parameter signed W23TO49 = 0;
parameter signed W23TO50 = 0;
parameter signed W23TO51 = 0;
parameter signed W23TO52 = 0;
parameter signed W23TO53 = 0;
parameter signed W23TO54 = 0;
parameter signed W23TO55 = 0;
parameter signed W23TO56 = 0;
parameter signed W23TO57 = 0;
parameter signed W23TO58 = 0;
parameter signed W23TO59 = 0;
parameter signed W23TO60 = 0;
parameter signed W23TO61 = 0;
parameter signed W23TO62 = 0;
parameter signed W23TO63 = 0;
parameter signed W24TO0 = 0;
parameter signed W24TO1 = 0;
parameter signed W24TO2 = 0;
parameter signed W24TO3 = 0;
parameter signed W24TO4 = 0;
parameter signed W24TO5 = 0;
parameter signed W24TO6 = 0;
parameter signed W24TO7 = 0;
parameter signed W24TO8 = 0;
parameter signed W24TO9 = 0;
parameter signed W24TO10 = 0;
parameter signed W24TO11 = 0;
parameter signed W24TO12 = 0;
parameter signed W24TO13 = 0;
parameter signed W24TO14 = 0;
parameter signed W24TO15 = 0;
parameter signed W24TO16 = 0;
parameter signed W24TO17 = 0;
parameter signed W24TO18 = 0;
parameter signed W24TO19 = 0;
parameter signed W24TO20 = 0;
parameter signed W24TO21 = 0;
parameter signed W24TO22 = 0;
parameter signed W24TO23 = 0;
parameter signed W24TO24 = 0;
parameter signed W24TO25 = 0;
parameter signed W24TO26 = 0;
parameter signed W24TO27 = 0;
parameter signed W24TO28 = 0;
parameter signed W24TO29 = 0;
parameter signed W24TO30 = 0;
parameter signed W24TO31 = 0;
parameter signed W24TO32 = 0;
parameter signed W24TO33 = 0;
parameter signed W24TO34 = 0;
parameter signed W24TO35 = 0;
parameter signed W24TO36 = 0;
parameter signed W24TO37 = 0;
parameter signed W24TO38 = 0;
parameter signed W24TO39 = 0;
parameter signed W24TO40 = 0;
parameter signed W24TO41 = 0;
parameter signed W24TO42 = 0;
parameter signed W24TO43 = 0;
parameter signed W24TO44 = 0;
parameter signed W24TO45 = 0;
parameter signed W24TO46 = 0;
parameter signed W24TO47 = 0;
parameter signed W24TO48 = 0;
parameter signed W24TO49 = 0;
parameter signed W24TO50 = 0;
parameter signed W24TO51 = 0;
parameter signed W24TO52 = 0;
parameter signed W24TO53 = 0;
parameter signed W24TO54 = 0;
parameter signed W24TO55 = 0;
parameter signed W24TO56 = 0;
parameter signed W24TO57 = 0;
parameter signed W24TO58 = 0;
parameter signed W24TO59 = 0;
parameter signed W24TO60 = 0;
parameter signed W24TO61 = 0;
parameter signed W24TO62 = 0;
parameter signed W24TO63 = 0;
parameter signed W25TO0 = 0;
parameter signed W25TO1 = 0;
parameter signed W25TO2 = 0;
parameter signed W25TO3 = 0;
parameter signed W25TO4 = 0;
parameter signed W25TO5 = 0;
parameter signed W25TO6 = 0;
parameter signed W25TO7 = 0;
parameter signed W25TO8 = 0;
parameter signed W25TO9 = 0;
parameter signed W25TO10 = 0;
parameter signed W25TO11 = 0;
parameter signed W25TO12 = 0;
parameter signed W25TO13 = 0;
parameter signed W25TO14 = 0;
parameter signed W25TO15 = 0;
parameter signed W25TO16 = 0;
parameter signed W25TO17 = 0;
parameter signed W25TO18 = 0;
parameter signed W25TO19 = 0;
parameter signed W25TO20 = 0;
parameter signed W25TO21 = 0;
parameter signed W25TO22 = 0;
parameter signed W25TO23 = 0;
parameter signed W25TO24 = 0;
parameter signed W25TO25 = 0;
parameter signed W25TO26 = 0;
parameter signed W25TO27 = 0;
parameter signed W25TO28 = 0;
parameter signed W25TO29 = 0;
parameter signed W25TO30 = 0;
parameter signed W25TO31 = 0;
parameter signed W25TO32 = 0;
parameter signed W25TO33 = 0;
parameter signed W25TO34 = 0;
parameter signed W25TO35 = 0;
parameter signed W25TO36 = 0;
parameter signed W25TO37 = 0;
parameter signed W25TO38 = 0;
parameter signed W25TO39 = 0;
parameter signed W25TO40 = 0;
parameter signed W25TO41 = 0;
parameter signed W25TO42 = 0;
parameter signed W25TO43 = 0;
parameter signed W25TO44 = 0;
parameter signed W25TO45 = 0;
parameter signed W25TO46 = 0;
parameter signed W25TO47 = 0;
parameter signed W25TO48 = 0;
parameter signed W25TO49 = 0;
parameter signed W25TO50 = 0;
parameter signed W25TO51 = 0;
parameter signed W25TO52 = 0;
parameter signed W25TO53 = 0;
parameter signed W25TO54 = 0;
parameter signed W25TO55 = 0;
parameter signed W25TO56 = 0;
parameter signed W25TO57 = 0;
parameter signed W25TO58 = 0;
parameter signed W25TO59 = 0;
parameter signed W25TO60 = 0;
parameter signed W25TO61 = 0;
parameter signed W25TO62 = 0;
parameter signed W25TO63 = 0;
parameter signed W26TO0 = 0;
parameter signed W26TO1 = 0;
parameter signed W26TO2 = 0;
parameter signed W26TO3 = 0;
parameter signed W26TO4 = 0;
parameter signed W26TO5 = 0;
parameter signed W26TO6 = 0;
parameter signed W26TO7 = 0;
parameter signed W26TO8 = 0;
parameter signed W26TO9 = 0;
parameter signed W26TO10 = 0;
parameter signed W26TO11 = 0;
parameter signed W26TO12 = 0;
parameter signed W26TO13 = 0;
parameter signed W26TO14 = 0;
parameter signed W26TO15 = 0;
parameter signed W26TO16 = 0;
parameter signed W26TO17 = 0;
parameter signed W26TO18 = 0;
parameter signed W26TO19 = 0;
parameter signed W26TO20 = 0;
parameter signed W26TO21 = 0;
parameter signed W26TO22 = 0;
parameter signed W26TO23 = 0;
parameter signed W26TO24 = 0;
parameter signed W26TO25 = 0;
parameter signed W26TO26 = 0;
parameter signed W26TO27 = 0;
parameter signed W26TO28 = 0;
parameter signed W26TO29 = 0;
parameter signed W26TO30 = 0;
parameter signed W26TO31 = 0;
parameter signed W26TO32 = 0;
parameter signed W26TO33 = 0;
parameter signed W26TO34 = 0;
parameter signed W26TO35 = 0;
parameter signed W26TO36 = 0;
parameter signed W26TO37 = 0;
parameter signed W26TO38 = 0;
parameter signed W26TO39 = 0;
parameter signed W26TO40 = 0;
parameter signed W26TO41 = 0;
parameter signed W26TO42 = 0;
parameter signed W26TO43 = 0;
parameter signed W26TO44 = 0;
parameter signed W26TO45 = 0;
parameter signed W26TO46 = 0;
parameter signed W26TO47 = 0;
parameter signed W26TO48 = 0;
parameter signed W26TO49 = 0;
parameter signed W26TO50 = 0;
parameter signed W26TO51 = 0;
parameter signed W26TO52 = 0;
parameter signed W26TO53 = 0;
parameter signed W26TO54 = 0;
parameter signed W26TO55 = 0;
parameter signed W26TO56 = 0;
parameter signed W26TO57 = 0;
parameter signed W26TO58 = 0;
parameter signed W26TO59 = 0;
parameter signed W26TO60 = 0;
parameter signed W26TO61 = 0;
parameter signed W26TO62 = 0;
parameter signed W26TO63 = 0;
parameter signed W27TO0 = 0;
parameter signed W27TO1 = 0;
parameter signed W27TO2 = 0;
parameter signed W27TO3 = 0;
parameter signed W27TO4 = 0;
parameter signed W27TO5 = 0;
parameter signed W27TO6 = 0;
parameter signed W27TO7 = 0;
parameter signed W27TO8 = 0;
parameter signed W27TO9 = 0;
parameter signed W27TO10 = 0;
parameter signed W27TO11 = 0;
parameter signed W27TO12 = 0;
parameter signed W27TO13 = 0;
parameter signed W27TO14 = 0;
parameter signed W27TO15 = 0;
parameter signed W27TO16 = 0;
parameter signed W27TO17 = 0;
parameter signed W27TO18 = 0;
parameter signed W27TO19 = 0;
parameter signed W27TO20 = 0;
parameter signed W27TO21 = 0;
parameter signed W27TO22 = 0;
parameter signed W27TO23 = 0;
parameter signed W27TO24 = 0;
parameter signed W27TO25 = 0;
parameter signed W27TO26 = 0;
parameter signed W27TO27 = 0;
parameter signed W27TO28 = 0;
parameter signed W27TO29 = 0;
parameter signed W27TO30 = 0;
parameter signed W27TO31 = 0;
parameter signed W27TO32 = 0;
parameter signed W27TO33 = 0;
parameter signed W27TO34 = 0;
parameter signed W27TO35 = 0;
parameter signed W27TO36 = 0;
parameter signed W27TO37 = 0;
parameter signed W27TO38 = 0;
parameter signed W27TO39 = 0;
parameter signed W27TO40 = 0;
parameter signed W27TO41 = 0;
parameter signed W27TO42 = 0;
parameter signed W27TO43 = 0;
parameter signed W27TO44 = 0;
parameter signed W27TO45 = 0;
parameter signed W27TO46 = 0;
parameter signed W27TO47 = 0;
parameter signed W27TO48 = 0;
parameter signed W27TO49 = 0;
parameter signed W27TO50 = 0;
parameter signed W27TO51 = 0;
parameter signed W27TO52 = 0;
parameter signed W27TO53 = 0;
parameter signed W27TO54 = 0;
parameter signed W27TO55 = 0;
parameter signed W27TO56 = 0;
parameter signed W27TO57 = 0;
parameter signed W27TO58 = 0;
parameter signed W27TO59 = 0;
parameter signed W27TO60 = 0;
parameter signed W27TO61 = 0;
parameter signed W27TO62 = 0;
parameter signed W27TO63 = 0;
parameter signed W28TO0 = 0;
parameter signed W28TO1 = 0;
parameter signed W28TO2 = 0;
parameter signed W28TO3 = 0;
parameter signed W28TO4 = 0;
parameter signed W28TO5 = 0;
parameter signed W28TO6 = 0;
parameter signed W28TO7 = 0;
parameter signed W28TO8 = 0;
parameter signed W28TO9 = 0;
parameter signed W28TO10 = 0;
parameter signed W28TO11 = 0;
parameter signed W28TO12 = 0;
parameter signed W28TO13 = 0;
parameter signed W28TO14 = 0;
parameter signed W28TO15 = 0;
parameter signed W28TO16 = 0;
parameter signed W28TO17 = 0;
parameter signed W28TO18 = 0;
parameter signed W28TO19 = 0;
parameter signed W28TO20 = 0;
parameter signed W28TO21 = 0;
parameter signed W28TO22 = 0;
parameter signed W28TO23 = 0;
parameter signed W28TO24 = 0;
parameter signed W28TO25 = 0;
parameter signed W28TO26 = 0;
parameter signed W28TO27 = 0;
parameter signed W28TO28 = 0;
parameter signed W28TO29 = 0;
parameter signed W28TO30 = 0;
parameter signed W28TO31 = 0;
parameter signed W28TO32 = 0;
parameter signed W28TO33 = 0;
parameter signed W28TO34 = 0;
parameter signed W28TO35 = 0;
parameter signed W28TO36 = 0;
parameter signed W28TO37 = 0;
parameter signed W28TO38 = 0;
parameter signed W28TO39 = 0;
parameter signed W28TO40 = 0;
parameter signed W28TO41 = 0;
parameter signed W28TO42 = 0;
parameter signed W28TO43 = 0;
parameter signed W28TO44 = 0;
parameter signed W28TO45 = 0;
parameter signed W28TO46 = 0;
parameter signed W28TO47 = 0;
parameter signed W28TO48 = 0;
parameter signed W28TO49 = 0;
parameter signed W28TO50 = 0;
parameter signed W28TO51 = 0;
parameter signed W28TO52 = 0;
parameter signed W28TO53 = 0;
parameter signed W28TO54 = 0;
parameter signed W28TO55 = 0;
parameter signed W28TO56 = 0;
parameter signed W28TO57 = 0;
parameter signed W28TO58 = 0;
parameter signed W28TO59 = 0;
parameter signed W28TO60 = 0;
parameter signed W28TO61 = 0;
parameter signed W28TO62 = 0;
parameter signed W28TO63 = 0;
parameter signed W29TO0 = 0;
parameter signed W29TO1 = 0;
parameter signed W29TO2 = 0;
parameter signed W29TO3 = 0;
parameter signed W29TO4 = 0;
parameter signed W29TO5 = 0;
parameter signed W29TO6 = 0;
parameter signed W29TO7 = 0;
parameter signed W29TO8 = 0;
parameter signed W29TO9 = 0;
parameter signed W29TO10 = 0;
parameter signed W29TO11 = 0;
parameter signed W29TO12 = 0;
parameter signed W29TO13 = 0;
parameter signed W29TO14 = 0;
parameter signed W29TO15 = 0;
parameter signed W29TO16 = 0;
parameter signed W29TO17 = 0;
parameter signed W29TO18 = 0;
parameter signed W29TO19 = 0;
parameter signed W29TO20 = 0;
parameter signed W29TO21 = 0;
parameter signed W29TO22 = 0;
parameter signed W29TO23 = 0;
parameter signed W29TO24 = 0;
parameter signed W29TO25 = 0;
parameter signed W29TO26 = 0;
parameter signed W29TO27 = 0;
parameter signed W29TO28 = 0;
parameter signed W29TO29 = 0;
parameter signed W29TO30 = 0;
parameter signed W29TO31 = 0;
parameter signed W29TO32 = 0;
parameter signed W29TO33 = 0;
parameter signed W29TO34 = 0;
parameter signed W29TO35 = 0;
parameter signed W29TO36 = 0;
parameter signed W29TO37 = 0;
parameter signed W29TO38 = 0;
parameter signed W29TO39 = 0;
parameter signed W29TO40 = 0;
parameter signed W29TO41 = 0;
parameter signed W29TO42 = 0;
parameter signed W29TO43 = 0;
parameter signed W29TO44 = 0;
parameter signed W29TO45 = 0;
parameter signed W29TO46 = 0;
parameter signed W29TO47 = 0;
parameter signed W29TO48 = 0;
parameter signed W29TO49 = 0;
parameter signed W29TO50 = 0;
parameter signed W29TO51 = 0;
parameter signed W29TO52 = 0;
parameter signed W29TO53 = 0;
parameter signed W29TO54 = 0;
parameter signed W29TO55 = 0;
parameter signed W29TO56 = 0;
parameter signed W29TO57 = 0;
parameter signed W29TO58 = 0;
parameter signed W29TO59 = 0;
parameter signed W29TO60 = 0;
parameter signed W29TO61 = 0;
parameter signed W29TO62 = 0;
parameter signed W29TO63 = 0;
parameter signed W30TO0 = 0;
parameter signed W30TO1 = 0;
parameter signed W30TO2 = 0;
parameter signed W30TO3 = 0;
parameter signed W30TO4 = 0;
parameter signed W30TO5 = 0;
parameter signed W30TO6 = 0;
parameter signed W30TO7 = 0;
parameter signed W30TO8 = 0;
parameter signed W30TO9 = 0;
parameter signed W30TO10 = 0;
parameter signed W30TO11 = 0;
parameter signed W30TO12 = 0;
parameter signed W30TO13 = 0;
parameter signed W30TO14 = 0;
parameter signed W30TO15 = 0;
parameter signed W30TO16 = 0;
parameter signed W30TO17 = 0;
parameter signed W30TO18 = 0;
parameter signed W30TO19 = 0;
parameter signed W30TO20 = 0;
parameter signed W30TO21 = 0;
parameter signed W30TO22 = 0;
parameter signed W30TO23 = 0;
parameter signed W30TO24 = 0;
parameter signed W30TO25 = 0;
parameter signed W30TO26 = 0;
parameter signed W30TO27 = 0;
parameter signed W30TO28 = 0;
parameter signed W30TO29 = 0;
parameter signed W30TO30 = 0;
parameter signed W30TO31 = 0;
parameter signed W30TO32 = 0;
parameter signed W30TO33 = 0;
parameter signed W30TO34 = 0;
parameter signed W30TO35 = 0;
parameter signed W30TO36 = 0;
parameter signed W30TO37 = 0;
parameter signed W30TO38 = 0;
parameter signed W30TO39 = 0;
parameter signed W30TO40 = 0;
parameter signed W30TO41 = 0;
parameter signed W30TO42 = 0;
parameter signed W30TO43 = 0;
parameter signed W30TO44 = 0;
parameter signed W30TO45 = 0;
parameter signed W30TO46 = 0;
parameter signed W30TO47 = 0;
parameter signed W30TO48 = 0;
parameter signed W30TO49 = 0;
parameter signed W30TO50 = 0;
parameter signed W30TO51 = 0;
parameter signed W30TO52 = 0;
parameter signed W30TO53 = 0;
parameter signed W30TO54 = 0;
parameter signed W30TO55 = 0;
parameter signed W30TO56 = 0;
parameter signed W30TO57 = 0;
parameter signed W30TO58 = 0;
parameter signed W30TO59 = 0;
parameter signed W30TO60 = 0;
parameter signed W30TO61 = 0;
parameter signed W30TO62 = 0;
parameter signed W30TO63 = 0;
parameter signed W31TO0 = 0;
parameter signed W31TO1 = 0;
parameter signed W31TO2 = 0;
parameter signed W31TO3 = 0;
parameter signed W31TO4 = 0;
parameter signed W31TO5 = 0;
parameter signed W31TO6 = 0;
parameter signed W31TO7 = 0;
parameter signed W31TO8 = 0;
parameter signed W31TO9 = 0;
parameter signed W31TO10 = 0;
parameter signed W31TO11 = 0;
parameter signed W31TO12 = 0;
parameter signed W31TO13 = 0;
parameter signed W31TO14 = 0;
parameter signed W31TO15 = 0;
parameter signed W31TO16 = 0;
parameter signed W31TO17 = 0;
parameter signed W31TO18 = 0;
parameter signed W31TO19 = 0;
parameter signed W31TO20 = 0;
parameter signed W31TO21 = 0;
parameter signed W31TO22 = 0;
parameter signed W31TO23 = 0;
parameter signed W31TO24 = 0;
parameter signed W31TO25 = 0;
parameter signed W31TO26 = 0;
parameter signed W31TO27 = 0;
parameter signed W31TO28 = 0;
parameter signed W31TO29 = 0;
parameter signed W31TO30 = 0;
parameter signed W31TO31 = 0;
parameter signed W31TO32 = 0;
parameter signed W31TO33 = 0;
parameter signed W31TO34 = 0;
parameter signed W31TO35 = 0;
parameter signed W31TO36 = 0;
parameter signed W31TO37 = 0;
parameter signed W31TO38 = 0;
parameter signed W31TO39 = 0;
parameter signed W31TO40 = 0;
parameter signed W31TO41 = 0;
parameter signed W31TO42 = 0;
parameter signed W31TO43 = 0;
parameter signed W31TO44 = 0;
parameter signed W31TO45 = 0;
parameter signed W31TO46 = 0;
parameter signed W31TO47 = 0;
parameter signed W31TO48 = 0;
parameter signed W31TO49 = 0;
parameter signed W31TO50 = 0;
parameter signed W31TO51 = 0;
parameter signed W31TO52 = 0;
parameter signed W31TO53 = 0;
parameter signed W31TO54 = 0;
parameter signed W31TO55 = 0;
parameter signed W31TO56 = 0;
parameter signed W31TO57 = 0;
parameter signed W31TO58 = 0;
parameter signed W31TO59 = 0;
parameter signed W31TO60 = 0;
parameter signed W31TO61 = 0;
parameter signed W31TO62 = 0;
parameter signed W31TO63 = 0;
parameter signed W32TO0 = 0;
parameter signed W32TO1 = 0;
parameter signed W32TO2 = 0;
parameter signed W32TO3 = 0;
parameter signed W32TO4 = 0;
parameter signed W32TO5 = 0;
parameter signed W32TO6 = 0;
parameter signed W32TO7 = 0;
parameter signed W32TO8 = 0;
parameter signed W32TO9 = 0;
parameter signed W32TO10 = 0;
parameter signed W32TO11 = 0;
parameter signed W32TO12 = 0;
parameter signed W32TO13 = 0;
parameter signed W32TO14 = 0;
parameter signed W32TO15 = 0;
parameter signed W32TO16 = 0;
parameter signed W32TO17 = 0;
parameter signed W32TO18 = 0;
parameter signed W32TO19 = 0;
parameter signed W32TO20 = 0;
parameter signed W32TO21 = 0;
parameter signed W32TO22 = 0;
parameter signed W32TO23 = 0;
parameter signed W32TO24 = 0;
parameter signed W32TO25 = 0;
parameter signed W32TO26 = 0;
parameter signed W32TO27 = 0;
parameter signed W32TO28 = 0;
parameter signed W32TO29 = 0;
parameter signed W32TO30 = 0;
parameter signed W32TO31 = 0;
parameter signed W32TO32 = 0;
parameter signed W32TO33 = 0;
parameter signed W32TO34 = 0;
parameter signed W32TO35 = 0;
parameter signed W32TO36 = 0;
parameter signed W32TO37 = 0;
parameter signed W32TO38 = 0;
parameter signed W32TO39 = 0;
parameter signed W32TO40 = 0;
parameter signed W32TO41 = 0;
parameter signed W32TO42 = 0;
parameter signed W32TO43 = 0;
parameter signed W32TO44 = 0;
parameter signed W32TO45 = 0;
parameter signed W32TO46 = 0;
parameter signed W32TO47 = 0;
parameter signed W32TO48 = 0;
parameter signed W32TO49 = 0;
parameter signed W32TO50 = 0;
parameter signed W32TO51 = 0;
parameter signed W32TO52 = 0;
parameter signed W32TO53 = 0;
parameter signed W32TO54 = 0;
parameter signed W32TO55 = 0;
parameter signed W32TO56 = 0;
parameter signed W32TO57 = 0;
parameter signed W32TO58 = 0;
parameter signed W32TO59 = 0;
parameter signed W32TO60 = 0;
parameter signed W32TO61 = 0;
parameter signed W32TO62 = 0;
parameter signed W32TO63 = 0;
parameter signed W33TO0 = 0;
parameter signed W33TO1 = 0;
parameter signed W33TO2 = 0;
parameter signed W33TO3 = 0;
parameter signed W33TO4 = 0;
parameter signed W33TO5 = 0;
parameter signed W33TO6 = 0;
parameter signed W33TO7 = 0;
parameter signed W33TO8 = 0;
parameter signed W33TO9 = 0;
parameter signed W33TO10 = 0;
parameter signed W33TO11 = 0;
parameter signed W33TO12 = 0;
parameter signed W33TO13 = 0;
parameter signed W33TO14 = 0;
parameter signed W33TO15 = 0;
parameter signed W33TO16 = 0;
parameter signed W33TO17 = 0;
parameter signed W33TO18 = 0;
parameter signed W33TO19 = 0;
parameter signed W33TO20 = 0;
parameter signed W33TO21 = 0;
parameter signed W33TO22 = 0;
parameter signed W33TO23 = 0;
parameter signed W33TO24 = 0;
parameter signed W33TO25 = 0;
parameter signed W33TO26 = 0;
parameter signed W33TO27 = 0;
parameter signed W33TO28 = 0;
parameter signed W33TO29 = 0;
parameter signed W33TO30 = 0;
parameter signed W33TO31 = 0;
parameter signed W33TO32 = 0;
parameter signed W33TO33 = 0;
parameter signed W33TO34 = 0;
parameter signed W33TO35 = 0;
parameter signed W33TO36 = 0;
parameter signed W33TO37 = 0;
parameter signed W33TO38 = 0;
parameter signed W33TO39 = 0;
parameter signed W33TO40 = 0;
parameter signed W33TO41 = 0;
parameter signed W33TO42 = 0;
parameter signed W33TO43 = 0;
parameter signed W33TO44 = 0;
parameter signed W33TO45 = 0;
parameter signed W33TO46 = 0;
parameter signed W33TO47 = 0;
parameter signed W33TO48 = 0;
parameter signed W33TO49 = 0;
parameter signed W33TO50 = 0;
parameter signed W33TO51 = 0;
parameter signed W33TO52 = 0;
parameter signed W33TO53 = 0;
parameter signed W33TO54 = 0;
parameter signed W33TO55 = 0;
parameter signed W33TO56 = 0;
parameter signed W33TO57 = 0;
parameter signed W33TO58 = 0;
parameter signed W33TO59 = 0;
parameter signed W33TO60 = 0;
parameter signed W33TO61 = 0;
parameter signed W33TO62 = 0;
parameter signed W33TO63 = 0;
parameter signed W34TO0 = 0;
parameter signed W34TO1 = 0;
parameter signed W34TO2 = 0;
parameter signed W34TO3 = 0;
parameter signed W34TO4 = 0;
parameter signed W34TO5 = 0;
parameter signed W34TO6 = 0;
parameter signed W34TO7 = 0;
parameter signed W34TO8 = 0;
parameter signed W34TO9 = 0;
parameter signed W34TO10 = 0;
parameter signed W34TO11 = 0;
parameter signed W34TO12 = 0;
parameter signed W34TO13 = 0;
parameter signed W34TO14 = 0;
parameter signed W34TO15 = 0;
parameter signed W34TO16 = 0;
parameter signed W34TO17 = 0;
parameter signed W34TO18 = 0;
parameter signed W34TO19 = 0;
parameter signed W34TO20 = 0;
parameter signed W34TO21 = 0;
parameter signed W34TO22 = 0;
parameter signed W34TO23 = 0;
parameter signed W34TO24 = 0;
parameter signed W34TO25 = 0;
parameter signed W34TO26 = 0;
parameter signed W34TO27 = 0;
parameter signed W34TO28 = 0;
parameter signed W34TO29 = 0;
parameter signed W34TO30 = 0;
parameter signed W34TO31 = 0;
parameter signed W34TO32 = 0;
parameter signed W34TO33 = 0;
parameter signed W34TO34 = 0;
parameter signed W34TO35 = 0;
parameter signed W34TO36 = 0;
parameter signed W34TO37 = 0;
parameter signed W34TO38 = 0;
parameter signed W34TO39 = 0;
parameter signed W34TO40 = 0;
parameter signed W34TO41 = 0;
parameter signed W34TO42 = 0;
parameter signed W34TO43 = 0;
parameter signed W34TO44 = 0;
parameter signed W34TO45 = 0;
parameter signed W34TO46 = 0;
parameter signed W34TO47 = 0;
parameter signed W34TO48 = 0;
parameter signed W34TO49 = 0;
parameter signed W34TO50 = 0;
parameter signed W34TO51 = 0;
parameter signed W34TO52 = 0;
parameter signed W34TO53 = 0;
parameter signed W34TO54 = 0;
parameter signed W34TO55 = 0;
parameter signed W34TO56 = 0;
parameter signed W34TO57 = 0;
parameter signed W34TO58 = 0;
parameter signed W34TO59 = 0;
parameter signed W34TO60 = 0;
parameter signed W34TO61 = 0;
parameter signed W34TO62 = 0;
parameter signed W34TO63 = 0;
parameter signed W35TO0 = 0;
parameter signed W35TO1 = 0;
parameter signed W35TO2 = 0;
parameter signed W35TO3 = 0;
parameter signed W35TO4 = 0;
parameter signed W35TO5 = 0;
parameter signed W35TO6 = 0;
parameter signed W35TO7 = 0;
parameter signed W35TO8 = 0;
parameter signed W35TO9 = 0;
parameter signed W35TO10 = 0;
parameter signed W35TO11 = 0;
parameter signed W35TO12 = 0;
parameter signed W35TO13 = 0;
parameter signed W35TO14 = 0;
parameter signed W35TO15 = 0;
parameter signed W35TO16 = 0;
parameter signed W35TO17 = 0;
parameter signed W35TO18 = 0;
parameter signed W35TO19 = 0;
parameter signed W35TO20 = 0;
parameter signed W35TO21 = 0;
parameter signed W35TO22 = 0;
parameter signed W35TO23 = 0;
parameter signed W35TO24 = 0;
parameter signed W35TO25 = 0;
parameter signed W35TO26 = 0;
parameter signed W35TO27 = 0;
parameter signed W35TO28 = 0;
parameter signed W35TO29 = 0;
parameter signed W35TO30 = 0;
parameter signed W35TO31 = 0;
parameter signed W35TO32 = 0;
parameter signed W35TO33 = 0;
parameter signed W35TO34 = 0;
parameter signed W35TO35 = 0;
parameter signed W35TO36 = 0;
parameter signed W35TO37 = 0;
parameter signed W35TO38 = 0;
parameter signed W35TO39 = 0;
parameter signed W35TO40 = 0;
parameter signed W35TO41 = 0;
parameter signed W35TO42 = 0;
parameter signed W35TO43 = 0;
parameter signed W35TO44 = 0;
parameter signed W35TO45 = 0;
parameter signed W35TO46 = 0;
parameter signed W35TO47 = 0;
parameter signed W35TO48 = 0;
parameter signed W35TO49 = 0;
parameter signed W35TO50 = 0;
parameter signed W35TO51 = 0;
parameter signed W35TO52 = 0;
parameter signed W35TO53 = 0;
parameter signed W35TO54 = 0;
parameter signed W35TO55 = 0;
parameter signed W35TO56 = 0;
parameter signed W35TO57 = 0;
parameter signed W35TO58 = 0;
parameter signed W35TO59 = 0;
parameter signed W35TO60 = 0;
parameter signed W35TO61 = 0;
parameter signed W35TO62 = 0;
parameter signed W35TO63 = 0;
parameter signed W36TO0 = 0;
parameter signed W36TO1 = 0;
parameter signed W36TO2 = 0;
parameter signed W36TO3 = 0;
parameter signed W36TO4 = 0;
parameter signed W36TO5 = 0;
parameter signed W36TO6 = 0;
parameter signed W36TO7 = 0;
parameter signed W36TO8 = 0;
parameter signed W36TO9 = 0;
parameter signed W36TO10 = 0;
parameter signed W36TO11 = 0;
parameter signed W36TO12 = 0;
parameter signed W36TO13 = 0;
parameter signed W36TO14 = 0;
parameter signed W36TO15 = 0;
parameter signed W36TO16 = 0;
parameter signed W36TO17 = 0;
parameter signed W36TO18 = 0;
parameter signed W36TO19 = 0;
parameter signed W36TO20 = 0;
parameter signed W36TO21 = 0;
parameter signed W36TO22 = 0;
parameter signed W36TO23 = 0;
parameter signed W36TO24 = 0;
parameter signed W36TO25 = 0;
parameter signed W36TO26 = 0;
parameter signed W36TO27 = 0;
parameter signed W36TO28 = 0;
parameter signed W36TO29 = 0;
parameter signed W36TO30 = 0;
parameter signed W36TO31 = 0;
parameter signed W36TO32 = 0;
parameter signed W36TO33 = 0;
parameter signed W36TO34 = 0;
parameter signed W36TO35 = 0;
parameter signed W36TO36 = 0;
parameter signed W36TO37 = 0;
parameter signed W36TO38 = 0;
parameter signed W36TO39 = 0;
parameter signed W36TO40 = 0;
parameter signed W36TO41 = 0;
parameter signed W36TO42 = 0;
parameter signed W36TO43 = 0;
parameter signed W36TO44 = 0;
parameter signed W36TO45 = 0;
parameter signed W36TO46 = 0;
parameter signed W36TO47 = 0;
parameter signed W36TO48 = 0;
parameter signed W36TO49 = 0;
parameter signed W36TO50 = 0;
parameter signed W36TO51 = 0;
parameter signed W36TO52 = 0;
parameter signed W36TO53 = 0;
parameter signed W36TO54 = 0;
parameter signed W36TO55 = 0;
parameter signed W36TO56 = 0;
parameter signed W36TO57 = 0;
parameter signed W36TO58 = 0;
parameter signed W36TO59 = 0;
parameter signed W36TO60 = 0;
parameter signed W36TO61 = 0;
parameter signed W36TO62 = 0;
parameter signed W36TO63 = 0;
parameter signed W37TO0 = 0;
parameter signed W37TO1 = 0;
parameter signed W37TO2 = 0;
parameter signed W37TO3 = 0;
parameter signed W37TO4 = 0;
parameter signed W37TO5 = 0;
parameter signed W37TO6 = 0;
parameter signed W37TO7 = 0;
parameter signed W37TO8 = 0;
parameter signed W37TO9 = 0;
parameter signed W37TO10 = 0;
parameter signed W37TO11 = 0;
parameter signed W37TO12 = 0;
parameter signed W37TO13 = 0;
parameter signed W37TO14 = 0;
parameter signed W37TO15 = 0;
parameter signed W37TO16 = 0;
parameter signed W37TO17 = 0;
parameter signed W37TO18 = 0;
parameter signed W37TO19 = 0;
parameter signed W37TO20 = 0;
parameter signed W37TO21 = 0;
parameter signed W37TO22 = 0;
parameter signed W37TO23 = 0;
parameter signed W37TO24 = 0;
parameter signed W37TO25 = 0;
parameter signed W37TO26 = 0;
parameter signed W37TO27 = 0;
parameter signed W37TO28 = 0;
parameter signed W37TO29 = 0;
parameter signed W37TO30 = 0;
parameter signed W37TO31 = 0;
parameter signed W37TO32 = 0;
parameter signed W37TO33 = 0;
parameter signed W37TO34 = 0;
parameter signed W37TO35 = 0;
parameter signed W37TO36 = 0;
parameter signed W37TO37 = 0;
parameter signed W37TO38 = 0;
parameter signed W37TO39 = 0;
parameter signed W37TO40 = 0;
parameter signed W37TO41 = 0;
parameter signed W37TO42 = 0;
parameter signed W37TO43 = 0;
parameter signed W37TO44 = 0;
parameter signed W37TO45 = 0;
parameter signed W37TO46 = 0;
parameter signed W37TO47 = 0;
parameter signed W37TO48 = 0;
parameter signed W37TO49 = 0;
parameter signed W37TO50 = 0;
parameter signed W37TO51 = 0;
parameter signed W37TO52 = 0;
parameter signed W37TO53 = 0;
parameter signed W37TO54 = 0;
parameter signed W37TO55 = 0;
parameter signed W37TO56 = 0;
parameter signed W37TO57 = 0;
parameter signed W37TO58 = 0;
parameter signed W37TO59 = 0;
parameter signed W37TO60 = 0;
parameter signed W37TO61 = 0;
parameter signed W37TO62 = 0;
parameter signed W37TO63 = 0;
parameter signed W38TO0 = 0;
parameter signed W38TO1 = 0;
parameter signed W38TO2 = 0;
parameter signed W38TO3 = 0;
parameter signed W38TO4 = 0;
parameter signed W38TO5 = 0;
parameter signed W38TO6 = 0;
parameter signed W38TO7 = 0;
parameter signed W38TO8 = 0;
parameter signed W38TO9 = 0;
parameter signed W38TO10 = 0;
parameter signed W38TO11 = 0;
parameter signed W38TO12 = 0;
parameter signed W38TO13 = 0;
parameter signed W38TO14 = 0;
parameter signed W38TO15 = 0;
parameter signed W38TO16 = 0;
parameter signed W38TO17 = 0;
parameter signed W38TO18 = 0;
parameter signed W38TO19 = 0;
parameter signed W38TO20 = 0;
parameter signed W38TO21 = 0;
parameter signed W38TO22 = 0;
parameter signed W38TO23 = 0;
parameter signed W38TO24 = 0;
parameter signed W38TO25 = 0;
parameter signed W38TO26 = 0;
parameter signed W38TO27 = 0;
parameter signed W38TO28 = 0;
parameter signed W38TO29 = 0;
parameter signed W38TO30 = 0;
parameter signed W38TO31 = 0;
parameter signed W38TO32 = 0;
parameter signed W38TO33 = 0;
parameter signed W38TO34 = 0;
parameter signed W38TO35 = 0;
parameter signed W38TO36 = 0;
parameter signed W38TO37 = 0;
parameter signed W38TO38 = 0;
parameter signed W38TO39 = 0;
parameter signed W38TO40 = 0;
parameter signed W38TO41 = 0;
parameter signed W38TO42 = 0;
parameter signed W38TO43 = 0;
parameter signed W38TO44 = 0;
parameter signed W38TO45 = 0;
parameter signed W38TO46 = 0;
parameter signed W38TO47 = 0;
parameter signed W38TO48 = 0;
parameter signed W38TO49 = 0;
parameter signed W38TO50 = 0;
parameter signed W38TO51 = 0;
parameter signed W38TO52 = 0;
parameter signed W38TO53 = 0;
parameter signed W38TO54 = 0;
parameter signed W38TO55 = 0;
parameter signed W38TO56 = 0;
parameter signed W38TO57 = 0;
parameter signed W38TO58 = 0;
parameter signed W38TO59 = 0;
parameter signed W38TO60 = 0;
parameter signed W38TO61 = 0;
parameter signed W38TO62 = 0;
parameter signed W38TO63 = 0;
parameter signed W39TO0 = 0;
parameter signed W39TO1 = 0;
parameter signed W39TO2 = 0;
parameter signed W39TO3 = 0;
parameter signed W39TO4 = 0;
parameter signed W39TO5 = 0;
parameter signed W39TO6 = 0;
parameter signed W39TO7 = 0;
parameter signed W39TO8 = 0;
parameter signed W39TO9 = 0;
parameter signed W39TO10 = 0;
parameter signed W39TO11 = 0;
parameter signed W39TO12 = 0;
parameter signed W39TO13 = 0;
parameter signed W39TO14 = 0;
parameter signed W39TO15 = 0;
parameter signed W39TO16 = 0;
parameter signed W39TO17 = 0;
parameter signed W39TO18 = 0;
parameter signed W39TO19 = 0;
parameter signed W39TO20 = 0;
parameter signed W39TO21 = 0;
parameter signed W39TO22 = 0;
parameter signed W39TO23 = 0;
parameter signed W39TO24 = 0;
parameter signed W39TO25 = 0;
parameter signed W39TO26 = 0;
parameter signed W39TO27 = 0;
parameter signed W39TO28 = 0;
parameter signed W39TO29 = 0;
parameter signed W39TO30 = 0;
parameter signed W39TO31 = 0;
parameter signed W39TO32 = 0;
parameter signed W39TO33 = 0;
parameter signed W39TO34 = 0;
parameter signed W39TO35 = 0;
parameter signed W39TO36 = 0;
parameter signed W39TO37 = 0;
parameter signed W39TO38 = 0;
parameter signed W39TO39 = 0;
parameter signed W39TO40 = 0;
parameter signed W39TO41 = 0;
parameter signed W39TO42 = 0;
parameter signed W39TO43 = 0;
parameter signed W39TO44 = 0;
parameter signed W39TO45 = 0;
parameter signed W39TO46 = 0;
parameter signed W39TO47 = 0;
parameter signed W39TO48 = 0;
parameter signed W39TO49 = 0;
parameter signed W39TO50 = 0;
parameter signed W39TO51 = 0;
parameter signed W39TO52 = 0;
parameter signed W39TO53 = 0;
parameter signed W39TO54 = 0;
parameter signed W39TO55 = 0;
parameter signed W39TO56 = 0;
parameter signed W39TO57 = 0;
parameter signed W39TO58 = 0;
parameter signed W39TO59 = 0;
parameter signed W39TO60 = 0;
parameter signed W39TO61 = 0;
parameter signed W39TO62 = 0;
parameter signed W39TO63 = 0;
parameter signed W40TO0 = 0;
parameter signed W40TO1 = 0;
parameter signed W40TO2 = 0;
parameter signed W40TO3 = 0;
parameter signed W40TO4 = 0;
parameter signed W40TO5 = 0;
parameter signed W40TO6 = 0;
parameter signed W40TO7 = 0;
parameter signed W40TO8 = 0;
parameter signed W40TO9 = 0;
parameter signed W40TO10 = 0;
parameter signed W40TO11 = 0;
parameter signed W40TO12 = 0;
parameter signed W40TO13 = 0;
parameter signed W40TO14 = 0;
parameter signed W40TO15 = 0;
parameter signed W40TO16 = 0;
parameter signed W40TO17 = 0;
parameter signed W40TO18 = 0;
parameter signed W40TO19 = 0;
parameter signed W40TO20 = 0;
parameter signed W40TO21 = 0;
parameter signed W40TO22 = 0;
parameter signed W40TO23 = 0;
parameter signed W40TO24 = 0;
parameter signed W40TO25 = 0;
parameter signed W40TO26 = 0;
parameter signed W40TO27 = 0;
parameter signed W40TO28 = 0;
parameter signed W40TO29 = 0;
parameter signed W40TO30 = 0;
parameter signed W40TO31 = 0;
parameter signed W40TO32 = 0;
parameter signed W40TO33 = 0;
parameter signed W40TO34 = 0;
parameter signed W40TO35 = 0;
parameter signed W40TO36 = 0;
parameter signed W40TO37 = 0;
parameter signed W40TO38 = 0;
parameter signed W40TO39 = 0;
parameter signed W40TO40 = 0;
parameter signed W40TO41 = 0;
parameter signed W40TO42 = 0;
parameter signed W40TO43 = 0;
parameter signed W40TO44 = 0;
parameter signed W40TO45 = 0;
parameter signed W40TO46 = 0;
parameter signed W40TO47 = 0;
parameter signed W40TO48 = 0;
parameter signed W40TO49 = 0;
parameter signed W40TO50 = 0;
parameter signed W40TO51 = 0;
parameter signed W40TO52 = 0;
parameter signed W40TO53 = 0;
parameter signed W40TO54 = 0;
parameter signed W40TO55 = 0;
parameter signed W40TO56 = 0;
parameter signed W40TO57 = 0;
parameter signed W40TO58 = 0;
parameter signed W40TO59 = 0;
parameter signed W40TO60 = 0;
parameter signed W40TO61 = 0;
parameter signed W40TO62 = 0;
parameter signed W40TO63 = 0;
parameter signed W41TO0 = 0;
parameter signed W41TO1 = 0;
parameter signed W41TO2 = 0;
parameter signed W41TO3 = 0;
parameter signed W41TO4 = 0;
parameter signed W41TO5 = 0;
parameter signed W41TO6 = 0;
parameter signed W41TO7 = 0;
parameter signed W41TO8 = 0;
parameter signed W41TO9 = 0;
parameter signed W41TO10 = 0;
parameter signed W41TO11 = 0;
parameter signed W41TO12 = 0;
parameter signed W41TO13 = 0;
parameter signed W41TO14 = 0;
parameter signed W41TO15 = 0;
parameter signed W41TO16 = 0;
parameter signed W41TO17 = 0;
parameter signed W41TO18 = 0;
parameter signed W41TO19 = 0;
parameter signed W41TO20 = 0;
parameter signed W41TO21 = 0;
parameter signed W41TO22 = 0;
parameter signed W41TO23 = 0;
parameter signed W41TO24 = 0;
parameter signed W41TO25 = 0;
parameter signed W41TO26 = 0;
parameter signed W41TO27 = 0;
parameter signed W41TO28 = 0;
parameter signed W41TO29 = 0;
parameter signed W41TO30 = 0;
parameter signed W41TO31 = 0;
parameter signed W41TO32 = 0;
parameter signed W41TO33 = 0;
parameter signed W41TO34 = 0;
parameter signed W41TO35 = 0;
parameter signed W41TO36 = 0;
parameter signed W41TO37 = 0;
parameter signed W41TO38 = 0;
parameter signed W41TO39 = 0;
parameter signed W41TO40 = 0;
parameter signed W41TO41 = 0;
parameter signed W41TO42 = 0;
parameter signed W41TO43 = 0;
parameter signed W41TO44 = 0;
parameter signed W41TO45 = 0;
parameter signed W41TO46 = 0;
parameter signed W41TO47 = 0;
parameter signed W41TO48 = 0;
parameter signed W41TO49 = 0;
parameter signed W41TO50 = 0;
parameter signed W41TO51 = 0;
parameter signed W41TO52 = 0;
parameter signed W41TO53 = 0;
parameter signed W41TO54 = 0;
parameter signed W41TO55 = 0;
parameter signed W41TO56 = 0;
parameter signed W41TO57 = 0;
parameter signed W41TO58 = 0;
parameter signed W41TO59 = 0;
parameter signed W41TO60 = 0;
parameter signed W41TO61 = 0;
parameter signed W41TO62 = 0;
parameter signed W41TO63 = 0;
parameter signed W42TO0 = 0;
parameter signed W42TO1 = 0;
parameter signed W42TO2 = 0;
parameter signed W42TO3 = 0;
parameter signed W42TO4 = 0;
parameter signed W42TO5 = 0;
parameter signed W42TO6 = 0;
parameter signed W42TO7 = 0;
parameter signed W42TO8 = 0;
parameter signed W42TO9 = 0;
parameter signed W42TO10 = 0;
parameter signed W42TO11 = 0;
parameter signed W42TO12 = 0;
parameter signed W42TO13 = 0;
parameter signed W42TO14 = 0;
parameter signed W42TO15 = 0;
parameter signed W42TO16 = 0;
parameter signed W42TO17 = 0;
parameter signed W42TO18 = 0;
parameter signed W42TO19 = 0;
parameter signed W42TO20 = 0;
parameter signed W42TO21 = 0;
parameter signed W42TO22 = 0;
parameter signed W42TO23 = 0;
parameter signed W42TO24 = 0;
parameter signed W42TO25 = 0;
parameter signed W42TO26 = 0;
parameter signed W42TO27 = 0;
parameter signed W42TO28 = 0;
parameter signed W42TO29 = 0;
parameter signed W42TO30 = 0;
parameter signed W42TO31 = 0;
parameter signed W42TO32 = 0;
parameter signed W42TO33 = 0;
parameter signed W42TO34 = 0;
parameter signed W42TO35 = 0;
parameter signed W42TO36 = 0;
parameter signed W42TO37 = 0;
parameter signed W42TO38 = 0;
parameter signed W42TO39 = 0;
parameter signed W42TO40 = 0;
parameter signed W42TO41 = 0;
parameter signed W42TO42 = 0;
parameter signed W42TO43 = 0;
parameter signed W42TO44 = 0;
parameter signed W42TO45 = 0;
parameter signed W42TO46 = 0;
parameter signed W42TO47 = 0;
parameter signed W42TO48 = 0;
parameter signed W42TO49 = 0;
parameter signed W42TO50 = 0;
parameter signed W42TO51 = 0;
parameter signed W42TO52 = 0;
parameter signed W42TO53 = 0;
parameter signed W42TO54 = 0;
parameter signed W42TO55 = 0;
parameter signed W42TO56 = 0;
parameter signed W42TO57 = 0;
parameter signed W42TO58 = 0;
parameter signed W42TO59 = 0;
parameter signed W42TO60 = 0;
parameter signed W42TO61 = 0;
parameter signed W42TO62 = 0;
parameter signed W42TO63 = 0;
parameter signed W43TO0 = 0;
parameter signed W43TO1 = 0;
parameter signed W43TO2 = 0;
parameter signed W43TO3 = 0;
parameter signed W43TO4 = 0;
parameter signed W43TO5 = 0;
parameter signed W43TO6 = 0;
parameter signed W43TO7 = 0;
parameter signed W43TO8 = 0;
parameter signed W43TO9 = 0;
parameter signed W43TO10 = 0;
parameter signed W43TO11 = 0;
parameter signed W43TO12 = 0;
parameter signed W43TO13 = 0;
parameter signed W43TO14 = 0;
parameter signed W43TO15 = 0;
parameter signed W43TO16 = 0;
parameter signed W43TO17 = 0;
parameter signed W43TO18 = 0;
parameter signed W43TO19 = 0;
parameter signed W43TO20 = 0;
parameter signed W43TO21 = 0;
parameter signed W43TO22 = 0;
parameter signed W43TO23 = 0;
parameter signed W43TO24 = 0;
parameter signed W43TO25 = 0;
parameter signed W43TO26 = 0;
parameter signed W43TO27 = 0;
parameter signed W43TO28 = 0;
parameter signed W43TO29 = 0;
parameter signed W43TO30 = 0;
parameter signed W43TO31 = 0;
parameter signed W43TO32 = 0;
parameter signed W43TO33 = 0;
parameter signed W43TO34 = 0;
parameter signed W43TO35 = 0;
parameter signed W43TO36 = 0;
parameter signed W43TO37 = 0;
parameter signed W43TO38 = 0;
parameter signed W43TO39 = 0;
parameter signed W43TO40 = 0;
parameter signed W43TO41 = 0;
parameter signed W43TO42 = 0;
parameter signed W43TO43 = 0;
parameter signed W43TO44 = 0;
parameter signed W43TO45 = 0;
parameter signed W43TO46 = 0;
parameter signed W43TO47 = 0;
parameter signed W43TO48 = 0;
parameter signed W43TO49 = 0;
parameter signed W43TO50 = 0;
parameter signed W43TO51 = 0;
parameter signed W43TO52 = 0;
parameter signed W43TO53 = 0;
parameter signed W43TO54 = 0;
parameter signed W43TO55 = 0;
parameter signed W43TO56 = 0;
parameter signed W43TO57 = 0;
parameter signed W43TO58 = 0;
parameter signed W43TO59 = 0;
parameter signed W43TO60 = 0;
parameter signed W43TO61 = 0;
parameter signed W43TO62 = 0;
parameter signed W43TO63 = 0;
parameter signed W44TO0 = 0;
parameter signed W44TO1 = 0;
parameter signed W44TO2 = 0;
parameter signed W44TO3 = 0;
parameter signed W44TO4 = 0;
parameter signed W44TO5 = 0;
parameter signed W44TO6 = 0;
parameter signed W44TO7 = 0;
parameter signed W44TO8 = 0;
parameter signed W44TO9 = 0;
parameter signed W44TO10 = 0;
parameter signed W44TO11 = 0;
parameter signed W44TO12 = 0;
parameter signed W44TO13 = 0;
parameter signed W44TO14 = 0;
parameter signed W44TO15 = 0;
parameter signed W44TO16 = 0;
parameter signed W44TO17 = 0;
parameter signed W44TO18 = 0;
parameter signed W44TO19 = 0;
parameter signed W44TO20 = 0;
parameter signed W44TO21 = 0;
parameter signed W44TO22 = 0;
parameter signed W44TO23 = 0;
parameter signed W44TO24 = 0;
parameter signed W44TO25 = 0;
parameter signed W44TO26 = 0;
parameter signed W44TO27 = 0;
parameter signed W44TO28 = 0;
parameter signed W44TO29 = 0;
parameter signed W44TO30 = 0;
parameter signed W44TO31 = 0;
parameter signed W44TO32 = 0;
parameter signed W44TO33 = 0;
parameter signed W44TO34 = 0;
parameter signed W44TO35 = 0;
parameter signed W44TO36 = 0;
parameter signed W44TO37 = 0;
parameter signed W44TO38 = 0;
parameter signed W44TO39 = 0;
parameter signed W44TO40 = 0;
parameter signed W44TO41 = 0;
parameter signed W44TO42 = 0;
parameter signed W44TO43 = 0;
parameter signed W44TO44 = 0;
parameter signed W44TO45 = 0;
parameter signed W44TO46 = 0;
parameter signed W44TO47 = 0;
parameter signed W44TO48 = 0;
parameter signed W44TO49 = 0;
parameter signed W44TO50 = 0;
parameter signed W44TO51 = 0;
parameter signed W44TO52 = 0;
parameter signed W44TO53 = 0;
parameter signed W44TO54 = 0;
parameter signed W44TO55 = 0;
parameter signed W44TO56 = 0;
parameter signed W44TO57 = 0;
parameter signed W44TO58 = 0;
parameter signed W44TO59 = 0;
parameter signed W44TO60 = 0;
parameter signed W44TO61 = 0;
parameter signed W44TO62 = 0;
parameter signed W44TO63 = 0;
parameter signed W45TO0 = 0;
parameter signed W45TO1 = 0;
parameter signed W45TO2 = 0;
parameter signed W45TO3 = 0;
parameter signed W45TO4 = 0;
parameter signed W45TO5 = 0;
parameter signed W45TO6 = 0;
parameter signed W45TO7 = 0;
parameter signed W45TO8 = 0;
parameter signed W45TO9 = 0;
parameter signed W45TO10 = 0;
parameter signed W45TO11 = 0;
parameter signed W45TO12 = 0;
parameter signed W45TO13 = 0;
parameter signed W45TO14 = 0;
parameter signed W45TO15 = 0;
parameter signed W45TO16 = 0;
parameter signed W45TO17 = 0;
parameter signed W45TO18 = 0;
parameter signed W45TO19 = 0;
parameter signed W45TO20 = 0;
parameter signed W45TO21 = 0;
parameter signed W45TO22 = 0;
parameter signed W45TO23 = 0;
parameter signed W45TO24 = 0;
parameter signed W45TO25 = 0;
parameter signed W45TO26 = 0;
parameter signed W45TO27 = 0;
parameter signed W45TO28 = 0;
parameter signed W45TO29 = 0;
parameter signed W45TO30 = 0;
parameter signed W45TO31 = 0;
parameter signed W45TO32 = 0;
parameter signed W45TO33 = 0;
parameter signed W45TO34 = 0;
parameter signed W45TO35 = 0;
parameter signed W45TO36 = 0;
parameter signed W45TO37 = 0;
parameter signed W45TO38 = 0;
parameter signed W45TO39 = 0;
parameter signed W45TO40 = 0;
parameter signed W45TO41 = 0;
parameter signed W45TO42 = 0;
parameter signed W45TO43 = 0;
parameter signed W45TO44 = 0;
parameter signed W45TO45 = 0;
parameter signed W45TO46 = 0;
parameter signed W45TO47 = 0;
parameter signed W45TO48 = 0;
parameter signed W45TO49 = 0;
parameter signed W45TO50 = 0;
parameter signed W45TO51 = 0;
parameter signed W45TO52 = 0;
parameter signed W45TO53 = 0;
parameter signed W45TO54 = 0;
parameter signed W45TO55 = 0;
parameter signed W45TO56 = 0;
parameter signed W45TO57 = 0;
parameter signed W45TO58 = 0;
parameter signed W45TO59 = 0;
parameter signed W45TO60 = 0;
parameter signed W45TO61 = 0;
parameter signed W45TO62 = 0;
parameter signed W45TO63 = 0;
parameter signed W46TO0 = 0;
parameter signed W46TO1 = 0;
parameter signed W46TO2 = 0;
parameter signed W46TO3 = 0;
parameter signed W46TO4 = 0;
parameter signed W46TO5 = 0;
parameter signed W46TO6 = 0;
parameter signed W46TO7 = 0;
parameter signed W46TO8 = 0;
parameter signed W46TO9 = 0;
parameter signed W46TO10 = 0;
parameter signed W46TO11 = 0;
parameter signed W46TO12 = 0;
parameter signed W46TO13 = 0;
parameter signed W46TO14 = 0;
parameter signed W46TO15 = 0;
parameter signed W46TO16 = 0;
parameter signed W46TO17 = 0;
parameter signed W46TO18 = 0;
parameter signed W46TO19 = 0;
parameter signed W46TO20 = 0;
parameter signed W46TO21 = 0;
parameter signed W46TO22 = 0;
parameter signed W46TO23 = 0;
parameter signed W46TO24 = 0;
parameter signed W46TO25 = 0;
parameter signed W46TO26 = 0;
parameter signed W46TO27 = 0;
parameter signed W46TO28 = 0;
parameter signed W46TO29 = 0;
parameter signed W46TO30 = 0;
parameter signed W46TO31 = 0;
parameter signed W46TO32 = 0;
parameter signed W46TO33 = 0;
parameter signed W46TO34 = 0;
parameter signed W46TO35 = 0;
parameter signed W46TO36 = 0;
parameter signed W46TO37 = 0;
parameter signed W46TO38 = 0;
parameter signed W46TO39 = 0;
parameter signed W46TO40 = 0;
parameter signed W46TO41 = 0;
parameter signed W46TO42 = 0;
parameter signed W46TO43 = 0;
parameter signed W46TO44 = 0;
parameter signed W46TO45 = 0;
parameter signed W46TO46 = 0;
parameter signed W46TO47 = 0;
parameter signed W46TO48 = 0;
parameter signed W46TO49 = 0;
parameter signed W46TO50 = 0;
parameter signed W46TO51 = 0;
parameter signed W46TO52 = 0;
parameter signed W46TO53 = 0;
parameter signed W46TO54 = 0;
parameter signed W46TO55 = 0;
parameter signed W46TO56 = 0;
parameter signed W46TO57 = 0;
parameter signed W46TO58 = 0;
parameter signed W46TO59 = 0;
parameter signed W46TO60 = 0;
parameter signed W46TO61 = 0;
parameter signed W46TO62 = 0;
parameter signed W46TO63 = 0;
parameter signed W47TO0 = 0;
parameter signed W47TO1 = 0;
parameter signed W47TO2 = 0;
parameter signed W47TO3 = 0;
parameter signed W47TO4 = 0;
parameter signed W47TO5 = 0;
parameter signed W47TO6 = 0;
parameter signed W47TO7 = 0;
parameter signed W47TO8 = 0;
parameter signed W47TO9 = 0;
parameter signed W47TO10 = 0;
parameter signed W47TO11 = 0;
parameter signed W47TO12 = 0;
parameter signed W47TO13 = 0;
parameter signed W47TO14 = 0;
parameter signed W47TO15 = 0;
parameter signed W47TO16 = 0;
parameter signed W47TO17 = 0;
parameter signed W47TO18 = 0;
parameter signed W47TO19 = 0;
parameter signed W47TO20 = 0;
parameter signed W47TO21 = 0;
parameter signed W47TO22 = 0;
parameter signed W47TO23 = 0;
parameter signed W47TO24 = 0;
parameter signed W47TO25 = 0;
parameter signed W47TO26 = 0;
parameter signed W47TO27 = 0;
parameter signed W47TO28 = 0;
parameter signed W47TO29 = 0;
parameter signed W47TO30 = 0;
parameter signed W47TO31 = 0;
parameter signed W47TO32 = 0;
parameter signed W47TO33 = 0;
parameter signed W47TO34 = 0;
parameter signed W47TO35 = 0;
parameter signed W47TO36 = 0;
parameter signed W47TO37 = 0;
parameter signed W47TO38 = 0;
parameter signed W47TO39 = 0;
parameter signed W47TO40 = 0;
parameter signed W47TO41 = 0;
parameter signed W47TO42 = 0;
parameter signed W47TO43 = 0;
parameter signed W47TO44 = 0;
parameter signed W47TO45 = 0;
parameter signed W47TO46 = 0;
parameter signed W47TO47 = 0;
parameter signed W47TO48 = 0;
parameter signed W47TO49 = 0;
parameter signed W47TO50 = 0;
parameter signed W47TO51 = 0;
parameter signed W47TO52 = 0;
parameter signed W47TO53 = 0;
parameter signed W47TO54 = 0;
parameter signed W47TO55 = 0;
parameter signed W47TO56 = 0;
parameter signed W47TO57 = 0;
parameter signed W47TO58 = 0;
parameter signed W47TO59 = 0;
parameter signed W47TO60 = 0;
parameter signed W47TO61 = 0;
parameter signed W47TO62 = 0;
parameter signed W47TO63 = 0;
parameter signed W48TO0 = 0;
parameter signed W48TO1 = 0;
parameter signed W48TO2 = 0;
parameter signed W48TO3 = 0;
parameter signed W48TO4 = 0;
parameter signed W48TO5 = 0;
parameter signed W48TO6 = 0;
parameter signed W48TO7 = 0;
parameter signed W48TO8 = 0;
parameter signed W48TO9 = 0;
parameter signed W48TO10 = 0;
parameter signed W48TO11 = 0;
parameter signed W48TO12 = 0;
parameter signed W48TO13 = 0;
parameter signed W48TO14 = 0;
parameter signed W48TO15 = 0;
parameter signed W48TO16 = 0;
parameter signed W48TO17 = 0;
parameter signed W48TO18 = 0;
parameter signed W48TO19 = 0;
parameter signed W48TO20 = 0;
parameter signed W48TO21 = 0;
parameter signed W48TO22 = 0;
parameter signed W48TO23 = 0;
parameter signed W48TO24 = 0;
parameter signed W48TO25 = 0;
parameter signed W48TO26 = 0;
parameter signed W48TO27 = 0;
parameter signed W48TO28 = 0;
parameter signed W48TO29 = 0;
parameter signed W48TO30 = 0;
parameter signed W48TO31 = 0;
parameter signed W48TO32 = 0;
parameter signed W48TO33 = 0;
parameter signed W48TO34 = 0;
parameter signed W48TO35 = 0;
parameter signed W48TO36 = 0;
parameter signed W48TO37 = 0;
parameter signed W48TO38 = 0;
parameter signed W48TO39 = 0;
parameter signed W48TO40 = 0;
parameter signed W48TO41 = 0;
parameter signed W48TO42 = 0;
parameter signed W48TO43 = 0;
parameter signed W48TO44 = 0;
parameter signed W48TO45 = 0;
parameter signed W48TO46 = 0;
parameter signed W48TO47 = 0;
parameter signed W48TO48 = 0;
parameter signed W48TO49 = 0;
parameter signed W48TO50 = 0;
parameter signed W48TO51 = 0;
parameter signed W48TO52 = 0;
parameter signed W48TO53 = 0;
parameter signed W48TO54 = 0;
parameter signed W48TO55 = 0;
parameter signed W48TO56 = 0;
parameter signed W48TO57 = 0;
parameter signed W48TO58 = 0;
parameter signed W48TO59 = 0;
parameter signed W48TO60 = 0;
parameter signed W48TO61 = 0;
parameter signed W48TO62 = 0;
parameter signed W48TO63 = 0;
parameter signed W49TO0 = 0;
parameter signed W49TO1 = 0;
parameter signed W49TO2 = 0;
parameter signed W49TO3 = 0;
parameter signed W49TO4 = 0;
parameter signed W49TO5 = 0;
parameter signed W49TO6 = 0;
parameter signed W49TO7 = 0;
parameter signed W49TO8 = 0;
parameter signed W49TO9 = 0;
parameter signed W49TO10 = 0;
parameter signed W49TO11 = 0;
parameter signed W49TO12 = 0;
parameter signed W49TO13 = 0;
parameter signed W49TO14 = 0;
parameter signed W49TO15 = 0;
parameter signed W49TO16 = 0;
parameter signed W49TO17 = 0;
parameter signed W49TO18 = 0;
parameter signed W49TO19 = 0;
parameter signed W49TO20 = 0;
parameter signed W49TO21 = 0;
parameter signed W49TO22 = 0;
parameter signed W49TO23 = 0;
parameter signed W49TO24 = 0;
parameter signed W49TO25 = 0;
parameter signed W49TO26 = 0;
parameter signed W49TO27 = 0;
parameter signed W49TO28 = 0;
parameter signed W49TO29 = 0;
parameter signed W49TO30 = 0;
parameter signed W49TO31 = 0;
parameter signed W49TO32 = 0;
parameter signed W49TO33 = 0;
parameter signed W49TO34 = 0;
parameter signed W49TO35 = 0;
parameter signed W49TO36 = 0;
parameter signed W49TO37 = 0;
parameter signed W49TO38 = 0;
parameter signed W49TO39 = 0;
parameter signed W49TO40 = 0;
parameter signed W49TO41 = 0;
parameter signed W49TO42 = 0;
parameter signed W49TO43 = 0;
parameter signed W49TO44 = 0;
parameter signed W49TO45 = 0;
parameter signed W49TO46 = 0;
parameter signed W49TO47 = 0;
parameter signed W49TO48 = 0;
parameter signed W49TO49 = 0;
parameter signed W49TO50 = 0;
parameter signed W49TO51 = 0;
parameter signed W49TO52 = 0;
parameter signed W49TO53 = 0;
parameter signed W49TO54 = 0;
parameter signed W49TO55 = 0;
parameter signed W49TO56 = 0;
parameter signed W49TO57 = 0;
parameter signed W49TO58 = 0;
parameter signed W49TO59 = 0;
parameter signed W49TO60 = 0;
parameter signed W49TO61 = 0;
parameter signed W49TO62 = 0;
parameter signed W49TO63 = 0;
parameter signed W50TO0 = 0;
parameter signed W50TO1 = 0;
parameter signed W50TO2 = 0;
parameter signed W50TO3 = 0;
parameter signed W50TO4 = 0;
parameter signed W50TO5 = 0;
parameter signed W50TO6 = 0;
parameter signed W50TO7 = 0;
parameter signed W50TO8 = 0;
parameter signed W50TO9 = 0;
parameter signed W50TO10 = 0;
parameter signed W50TO11 = 0;
parameter signed W50TO12 = 0;
parameter signed W50TO13 = 0;
parameter signed W50TO14 = 0;
parameter signed W50TO15 = 0;
parameter signed W50TO16 = 0;
parameter signed W50TO17 = 0;
parameter signed W50TO18 = 0;
parameter signed W50TO19 = 0;
parameter signed W50TO20 = 0;
parameter signed W50TO21 = 0;
parameter signed W50TO22 = 0;
parameter signed W50TO23 = 0;
parameter signed W50TO24 = 0;
parameter signed W50TO25 = 0;
parameter signed W50TO26 = 0;
parameter signed W50TO27 = 0;
parameter signed W50TO28 = 0;
parameter signed W50TO29 = 0;
parameter signed W50TO30 = 0;
parameter signed W50TO31 = 0;
parameter signed W50TO32 = 0;
parameter signed W50TO33 = 0;
parameter signed W50TO34 = 0;
parameter signed W50TO35 = 0;
parameter signed W50TO36 = 0;
parameter signed W50TO37 = 0;
parameter signed W50TO38 = 0;
parameter signed W50TO39 = 0;
parameter signed W50TO40 = 0;
parameter signed W50TO41 = 0;
parameter signed W50TO42 = 0;
parameter signed W50TO43 = 0;
parameter signed W50TO44 = 0;
parameter signed W50TO45 = 0;
parameter signed W50TO46 = 0;
parameter signed W50TO47 = 0;
parameter signed W50TO48 = 0;
parameter signed W50TO49 = 0;
parameter signed W50TO50 = 0;
parameter signed W50TO51 = 0;
parameter signed W50TO52 = 0;
parameter signed W50TO53 = 0;
parameter signed W50TO54 = 0;
parameter signed W50TO55 = 0;
parameter signed W50TO56 = 0;
parameter signed W50TO57 = 0;
parameter signed W50TO58 = 0;
parameter signed W50TO59 = 0;
parameter signed W50TO60 = 0;
parameter signed W50TO61 = 0;
parameter signed W50TO62 = 0;
parameter signed W50TO63 = 0;
parameter signed W51TO0 = 0;
parameter signed W51TO1 = 0;
parameter signed W51TO2 = 0;
parameter signed W51TO3 = 0;
parameter signed W51TO4 = 0;
parameter signed W51TO5 = 0;
parameter signed W51TO6 = 0;
parameter signed W51TO7 = 0;
parameter signed W51TO8 = 0;
parameter signed W51TO9 = 0;
parameter signed W51TO10 = 0;
parameter signed W51TO11 = 0;
parameter signed W51TO12 = 0;
parameter signed W51TO13 = 0;
parameter signed W51TO14 = 0;
parameter signed W51TO15 = 0;
parameter signed W51TO16 = 0;
parameter signed W51TO17 = 0;
parameter signed W51TO18 = 0;
parameter signed W51TO19 = 0;
parameter signed W51TO20 = 0;
parameter signed W51TO21 = 0;
parameter signed W51TO22 = 0;
parameter signed W51TO23 = 0;
parameter signed W51TO24 = 0;
parameter signed W51TO25 = 0;
parameter signed W51TO26 = 0;
parameter signed W51TO27 = 0;
parameter signed W51TO28 = 0;
parameter signed W51TO29 = 0;
parameter signed W51TO30 = 0;
parameter signed W51TO31 = 0;
parameter signed W51TO32 = 0;
parameter signed W51TO33 = 0;
parameter signed W51TO34 = 0;
parameter signed W51TO35 = 0;
parameter signed W51TO36 = 0;
parameter signed W51TO37 = 0;
parameter signed W51TO38 = 0;
parameter signed W51TO39 = 0;
parameter signed W51TO40 = 0;
parameter signed W51TO41 = 0;
parameter signed W51TO42 = 0;
parameter signed W51TO43 = 0;
parameter signed W51TO44 = 0;
parameter signed W51TO45 = 0;
parameter signed W51TO46 = 0;
parameter signed W51TO47 = 0;
parameter signed W51TO48 = 0;
parameter signed W51TO49 = 0;
parameter signed W51TO50 = 0;
parameter signed W51TO51 = 0;
parameter signed W51TO52 = 0;
parameter signed W51TO53 = 0;
parameter signed W51TO54 = 0;
parameter signed W51TO55 = 0;
parameter signed W51TO56 = 0;
parameter signed W51TO57 = 0;
parameter signed W51TO58 = 0;
parameter signed W51TO59 = 0;
parameter signed W51TO60 = 0;
parameter signed W51TO61 = 0;
parameter signed W51TO62 = 0;
parameter signed W51TO63 = 0;
parameter signed W52TO0 = 0;
parameter signed W52TO1 = 0;
parameter signed W52TO2 = 0;
parameter signed W52TO3 = 0;
parameter signed W52TO4 = 0;
parameter signed W52TO5 = 0;
parameter signed W52TO6 = 0;
parameter signed W52TO7 = 0;
parameter signed W52TO8 = 0;
parameter signed W52TO9 = 0;
parameter signed W52TO10 = 0;
parameter signed W52TO11 = 0;
parameter signed W52TO12 = 0;
parameter signed W52TO13 = 0;
parameter signed W52TO14 = 0;
parameter signed W52TO15 = 0;
parameter signed W52TO16 = 0;
parameter signed W52TO17 = 0;
parameter signed W52TO18 = 0;
parameter signed W52TO19 = 0;
parameter signed W52TO20 = 0;
parameter signed W52TO21 = 0;
parameter signed W52TO22 = 0;
parameter signed W52TO23 = 0;
parameter signed W52TO24 = 0;
parameter signed W52TO25 = 0;
parameter signed W52TO26 = 0;
parameter signed W52TO27 = 0;
parameter signed W52TO28 = 0;
parameter signed W52TO29 = 0;
parameter signed W52TO30 = 0;
parameter signed W52TO31 = 0;
parameter signed W52TO32 = 0;
parameter signed W52TO33 = 0;
parameter signed W52TO34 = 0;
parameter signed W52TO35 = 0;
parameter signed W52TO36 = 0;
parameter signed W52TO37 = 0;
parameter signed W52TO38 = 0;
parameter signed W52TO39 = 0;
parameter signed W52TO40 = 0;
parameter signed W52TO41 = 0;
parameter signed W52TO42 = 0;
parameter signed W52TO43 = 0;
parameter signed W52TO44 = 0;
parameter signed W52TO45 = 0;
parameter signed W52TO46 = 0;
parameter signed W52TO47 = 0;
parameter signed W52TO48 = 0;
parameter signed W52TO49 = 0;
parameter signed W52TO50 = 0;
parameter signed W52TO51 = 0;
parameter signed W52TO52 = 0;
parameter signed W52TO53 = 0;
parameter signed W52TO54 = 0;
parameter signed W52TO55 = 0;
parameter signed W52TO56 = 0;
parameter signed W52TO57 = 0;
parameter signed W52TO58 = 0;
parameter signed W52TO59 = 0;
parameter signed W52TO60 = 0;
parameter signed W52TO61 = 0;
parameter signed W52TO62 = 0;
parameter signed W52TO63 = 0;
parameter signed W53TO0 = 0;
parameter signed W53TO1 = 0;
parameter signed W53TO2 = 0;
parameter signed W53TO3 = 0;
parameter signed W53TO4 = 0;
parameter signed W53TO5 = 0;
parameter signed W53TO6 = 0;
parameter signed W53TO7 = 0;
parameter signed W53TO8 = 0;
parameter signed W53TO9 = 0;
parameter signed W53TO10 = 0;
parameter signed W53TO11 = 0;
parameter signed W53TO12 = 0;
parameter signed W53TO13 = 0;
parameter signed W53TO14 = 0;
parameter signed W53TO15 = 0;
parameter signed W53TO16 = 0;
parameter signed W53TO17 = 0;
parameter signed W53TO18 = 0;
parameter signed W53TO19 = 0;
parameter signed W53TO20 = 0;
parameter signed W53TO21 = 0;
parameter signed W53TO22 = 0;
parameter signed W53TO23 = 0;
parameter signed W53TO24 = 0;
parameter signed W53TO25 = 0;
parameter signed W53TO26 = 0;
parameter signed W53TO27 = 0;
parameter signed W53TO28 = 0;
parameter signed W53TO29 = 0;
parameter signed W53TO30 = 0;
parameter signed W53TO31 = 0;
parameter signed W53TO32 = 0;
parameter signed W53TO33 = 0;
parameter signed W53TO34 = 0;
parameter signed W53TO35 = 0;
parameter signed W53TO36 = 0;
parameter signed W53TO37 = 0;
parameter signed W53TO38 = 0;
parameter signed W53TO39 = 0;
parameter signed W53TO40 = 0;
parameter signed W53TO41 = 0;
parameter signed W53TO42 = 0;
parameter signed W53TO43 = 0;
parameter signed W53TO44 = 0;
parameter signed W53TO45 = 0;
parameter signed W53TO46 = 0;
parameter signed W53TO47 = 0;
parameter signed W53TO48 = 0;
parameter signed W53TO49 = 0;
parameter signed W53TO50 = 0;
parameter signed W53TO51 = 0;
parameter signed W53TO52 = 0;
parameter signed W53TO53 = 0;
parameter signed W53TO54 = 0;
parameter signed W53TO55 = 0;
parameter signed W53TO56 = 0;
parameter signed W53TO57 = 0;
parameter signed W53TO58 = 0;
parameter signed W53TO59 = 0;
parameter signed W53TO60 = 0;
parameter signed W53TO61 = 0;
parameter signed W53TO62 = 0;
parameter signed W53TO63 = 0;
parameter signed W54TO0 = 0;
parameter signed W54TO1 = 0;
parameter signed W54TO2 = 0;
parameter signed W54TO3 = 0;
parameter signed W54TO4 = 0;
parameter signed W54TO5 = 0;
parameter signed W54TO6 = 0;
parameter signed W54TO7 = 0;
parameter signed W54TO8 = 0;
parameter signed W54TO9 = 0;
parameter signed W54TO10 = 0;
parameter signed W54TO11 = 0;
parameter signed W54TO12 = 0;
parameter signed W54TO13 = 0;
parameter signed W54TO14 = 0;
parameter signed W54TO15 = 0;
parameter signed W54TO16 = 0;
parameter signed W54TO17 = 0;
parameter signed W54TO18 = 0;
parameter signed W54TO19 = 0;
parameter signed W54TO20 = 0;
parameter signed W54TO21 = 0;
parameter signed W54TO22 = 0;
parameter signed W54TO23 = 0;
parameter signed W54TO24 = 0;
parameter signed W54TO25 = 0;
parameter signed W54TO26 = 0;
parameter signed W54TO27 = 0;
parameter signed W54TO28 = 0;
parameter signed W54TO29 = 0;
parameter signed W54TO30 = 0;
parameter signed W54TO31 = 0;
parameter signed W54TO32 = 0;
parameter signed W54TO33 = 0;
parameter signed W54TO34 = 0;
parameter signed W54TO35 = 0;
parameter signed W54TO36 = 0;
parameter signed W54TO37 = 0;
parameter signed W54TO38 = 0;
parameter signed W54TO39 = 0;
parameter signed W54TO40 = 0;
parameter signed W54TO41 = 0;
parameter signed W54TO42 = 0;
parameter signed W54TO43 = 0;
parameter signed W54TO44 = 0;
parameter signed W54TO45 = 0;
parameter signed W54TO46 = 0;
parameter signed W54TO47 = 0;
parameter signed W54TO48 = 0;
parameter signed W54TO49 = 0;
parameter signed W54TO50 = 0;
parameter signed W54TO51 = 0;
parameter signed W54TO52 = 0;
parameter signed W54TO53 = 0;
parameter signed W54TO54 = 0;
parameter signed W54TO55 = 0;
parameter signed W54TO56 = 0;
parameter signed W54TO57 = 0;
parameter signed W54TO58 = 0;
parameter signed W54TO59 = 0;
parameter signed W54TO60 = 0;
parameter signed W54TO61 = 0;
parameter signed W54TO62 = 0;
parameter signed W54TO63 = 0;
parameter signed W55TO0 = 0;
parameter signed W55TO1 = 0;
parameter signed W55TO2 = 0;
parameter signed W55TO3 = 0;
parameter signed W55TO4 = 0;
parameter signed W55TO5 = 0;
parameter signed W55TO6 = 0;
parameter signed W55TO7 = 0;
parameter signed W55TO8 = 0;
parameter signed W55TO9 = 0;
parameter signed W55TO10 = 0;
parameter signed W55TO11 = 0;
parameter signed W55TO12 = 0;
parameter signed W55TO13 = 0;
parameter signed W55TO14 = 0;
parameter signed W55TO15 = 0;
parameter signed W55TO16 = 0;
parameter signed W55TO17 = 0;
parameter signed W55TO18 = 0;
parameter signed W55TO19 = 0;
parameter signed W55TO20 = 0;
parameter signed W55TO21 = 0;
parameter signed W55TO22 = 0;
parameter signed W55TO23 = 0;
parameter signed W55TO24 = 0;
parameter signed W55TO25 = 0;
parameter signed W55TO26 = 0;
parameter signed W55TO27 = 0;
parameter signed W55TO28 = 0;
parameter signed W55TO29 = 0;
parameter signed W55TO30 = 0;
parameter signed W55TO31 = 0;
parameter signed W55TO32 = 0;
parameter signed W55TO33 = 0;
parameter signed W55TO34 = 0;
parameter signed W55TO35 = 0;
parameter signed W55TO36 = 0;
parameter signed W55TO37 = 0;
parameter signed W55TO38 = 0;
parameter signed W55TO39 = 0;
parameter signed W55TO40 = 0;
parameter signed W55TO41 = 0;
parameter signed W55TO42 = 0;
parameter signed W55TO43 = 0;
parameter signed W55TO44 = 0;
parameter signed W55TO45 = 0;
parameter signed W55TO46 = 0;
parameter signed W55TO47 = 0;
parameter signed W55TO48 = 0;
parameter signed W55TO49 = 0;
parameter signed W55TO50 = 0;
parameter signed W55TO51 = 0;
parameter signed W55TO52 = 0;
parameter signed W55TO53 = 0;
parameter signed W55TO54 = 0;
parameter signed W55TO55 = 0;
parameter signed W55TO56 = 0;
parameter signed W55TO57 = 0;
parameter signed W55TO58 = 0;
parameter signed W55TO59 = 0;
parameter signed W55TO60 = 0;
parameter signed W55TO61 = 0;
parameter signed W55TO62 = 0;
parameter signed W55TO63 = 0;
parameter signed W56TO0 = 0;
parameter signed W56TO1 = 0;
parameter signed W56TO2 = 0;
parameter signed W56TO3 = 0;
parameter signed W56TO4 = 0;
parameter signed W56TO5 = 0;
parameter signed W56TO6 = 0;
parameter signed W56TO7 = 0;
parameter signed W56TO8 = 0;
parameter signed W56TO9 = 0;
parameter signed W56TO10 = 0;
parameter signed W56TO11 = 0;
parameter signed W56TO12 = 0;
parameter signed W56TO13 = 0;
parameter signed W56TO14 = 0;
parameter signed W56TO15 = 0;
parameter signed W56TO16 = 0;
parameter signed W56TO17 = 0;
parameter signed W56TO18 = 0;
parameter signed W56TO19 = 0;
parameter signed W56TO20 = 0;
parameter signed W56TO21 = 0;
parameter signed W56TO22 = 0;
parameter signed W56TO23 = 0;
parameter signed W56TO24 = 0;
parameter signed W56TO25 = 0;
parameter signed W56TO26 = 0;
parameter signed W56TO27 = 0;
parameter signed W56TO28 = 0;
parameter signed W56TO29 = 0;
parameter signed W56TO30 = 0;
parameter signed W56TO31 = 0;
parameter signed W56TO32 = 0;
parameter signed W56TO33 = 0;
parameter signed W56TO34 = 0;
parameter signed W56TO35 = 0;
parameter signed W56TO36 = 0;
parameter signed W56TO37 = 0;
parameter signed W56TO38 = 0;
parameter signed W56TO39 = 0;
parameter signed W56TO40 = 0;
parameter signed W56TO41 = 0;
parameter signed W56TO42 = 0;
parameter signed W56TO43 = 0;
parameter signed W56TO44 = 0;
parameter signed W56TO45 = 0;
parameter signed W56TO46 = 0;
parameter signed W56TO47 = 0;
parameter signed W56TO48 = 0;
parameter signed W56TO49 = 0;
parameter signed W56TO50 = 0;
parameter signed W56TO51 = 0;
parameter signed W56TO52 = 0;
parameter signed W56TO53 = 0;
parameter signed W56TO54 = 0;
parameter signed W56TO55 = 0;
parameter signed W56TO56 = 0;
parameter signed W56TO57 = 0;
parameter signed W56TO58 = 0;
parameter signed W56TO59 = 0;
parameter signed W56TO60 = 0;
parameter signed W56TO61 = 0;
parameter signed W56TO62 = 0;
parameter signed W56TO63 = 0;
parameter signed W57TO0 = 0;
parameter signed W57TO1 = 0;
parameter signed W57TO2 = 0;
parameter signed W57TO3 = 0;
parameter signed W57TO4 = 0;
parameter signed W57TO5 = 0;
parameter signed W57TO6 = 0;
parameter signed W57TO7 = 0;
parameter signed W57TO8 = 0;
parameter signed W57TO9 = 0;
parameter signed W57TO10 = 0;
parameter signed W57TO11 = 0;
parameter signed W57TO12 = 0;
parameter signed W57TO13 = 0;
parameter signed W57TO14 = 0;
parameter signed W57TO15 = 0;
parameter signed W57TO16 = 0;
parameter signed W57TO17 = 0;
parameter signed W57TO18 = 0;
parameter signed W57TO19 = 0;
parameter signed W57TO20 = 0;
parameter signed W57TO21 = 0;
parameter signed W57TO22 = 0;
parameter signed W57TO23 = 0;
parameter signed W57TO24 = 0;
parameter signed W57TO25 = 0;
parameter signed W57TO26 = 0;
parameter signed W57TO27 = 0;
parameter signed W57TO28 = 0;
parameter signed W57TO29 = 0;
parameter signed W57TO30 = 0;
parameter signed W57TO31 = 0;
parameter signed W57TO32 = 0;
parameter signed W57TO33 = 0;
parameter signed W57TO34 = 0;
parameter signed W57TO35 = 0;
parameter signed W57TO36 = 0;
parameter signed W57TO37 = 0;
parameter signed W57TO38 = 0;
parameter signed W57TO39 = 0;
parameter signed W57TO40 = 0;
parameter signed W57TO41 = 0;
parameter signed W57TO42 = 0;
parameter signed W57TO43 = 0;
parameter signed W57TO44 = 0;
parameter signed W57TO45 = 0;
parameter signed W57TO46 = 0;
parameter signed W57TO47 = 0;
parameter signed W57TO48 = 0;
parameter signed W57TO49 = 0;
parameter signed W57TO50 = 0;
parameter signed W57TO51 = 0;
parameter signed W57TO52 = 0;
parameter signed W57TO53 = 0;
parameter signed W57TO54 = 0;
parameter signed W57TO55 = 0;
parameter signed W57TO56 = 0;
parameter signed W57TO57 = 0;
parameter signed W57TO58 = 0;
parameter signed W57TO59 = 0;
parameter signed W57TO60 = 0;
parameter signed W57TO61 = 0;
parameter signed W57TO62 = 0;
parameter signed W57TO63 = 0;
parameter signed W58TO0 = 0;
parameter signed W58TO1 = 0;
parameter signed W58TO2 = 0;
parameter signed W58TO3 = 0;
parameter signed W58TO4 = 0;
parameter signed W58TO5 = 0;
parameter signed W58TO6 = 0;
parameter signed W58TO7 = 0;
parameter signed W58TO8 = 0;
parameter signed W58TO9 = 0;
parameter signed W58TO10 = 0;
parameter signed W58TO11 = 0;
parameter signed W58TO12 = 0;
parameter signed W58TO13 = 0;
parameter signed W58TO14 = 0;
parameter signed W58TO15 = 0;
parameter signed W58TO16 = 0;
parameter signed W58TO17 = 0;
parameter signed W58TO18 = 0;
parameter signed W58TO19 = 0;
parameter signed W58TO20 = 0;
parameter signed W58TO21 = 0;
parameter signed W58TO22 = 0;
parameter signed W58TO23 = 0;
parameter signed W58TO24 = 0;
parameter signed W58TO25 = 0;
parameter signed W58TO26 = 0;
parameter signed W58TO27 = 0;
parameter signed W58TO28 = 0;
parameter signed W58TO29 = 0;
parameter signed W58TO30 = 0;
parameter signed W58TO31 = 0;
parameter signed W58TO32 = 0;
parameter signed W58TO33 = 0;
parameter signed W58TO34 = 0;
parameter signed W58TO35 = 0;
parameter signed W58TO36 = 0;
parameter signed W58TO37 = 0;
parameter signed W58TO38 = 0;
parameter signed W58TO39 = 0;
parameter signed W58TO40 = 0;
parameter signed W58TO41 = 0;
parameter signed W58TO42 = 0;
parameter signed W58TO43 = 0;
parameter signed W58TO44 = 0;
parameter signed W58TO45 = 0;
parameter signed W58TO46 = 0;
parameter signed W58TO47 = 0;
parameter signed W58TO48 = 0;
parameter signed W58TO49 = 0;
parameter signed W58TO50 = 0;
parameter signed W58TO51 = 0;
parameter signed W58TO52 = 0;
parameter signed W58TO53 = 0;
parameter signed W58TO54 = 0;
parameter signed W58TO55 = 0;
parameter signed W58TO56 = 0;
parameter signed W58TO57 = 0;
parameter signed W58TO58 = 0;
parameter signed W58TO59 = 0;
parameter signed W58TO60 = 0;
parameter signed W58TO61 = 0;
parameter signed W58TO62 = 0;
parameter signed W58TO63 = 0;
parameter signed W59TO0 = 0;
parameter signed W59TO1 = 0;
parameter signed W59TO2 = 0;
parameter signed W59TO3 = 0;
parameter signed W59TO4 = 0;
parameter signed W59TO5 = 0;
parameter signed W59TO6 = 0;
parameter signed W59TO7 = 0;
parameter signed W59TO8 = 0;
parameter signed W59TO9 = 0;
parameter signed W59TO10 = 0;
parameter signed W59TO11 = 0;
parameter signed W59TO12 = 0;
parameter signed W59TO13 = 0;
parameter signed W59TO14 = 0;
parameter signed W59TO15 = 0;
parameter signed W59TO16 = 0;
parameter signed W59TO17 = 0;
parameter signed W59TO18 = 0;
parameter signed W59TO19 = 0;
parameter signed W59TO20 = 0;
parameter signed W59TO21 = 0;
parameter signed W59TO22 = 0;
parameter signed W59TO23 = 0;
parameter signed W59TO24 = 0;
parameter signed W59TO25 = 0;
parameter signed W59TO26 = 0;
parameter signed W59TO27 = 0;
parameter signed W59TO28 = 0;
parameter signed W59TO29 = 0;
parameter signed W59TO30 = 0;
parameter signed W59TO31 = 0;
parameter signed W59TO32 = 0;
parameter signed W59TO33 = 0;
parameter signed W59TO34 = 0;
parameter signed W59TO35 = 0;
parameter signed W59TO36 = 0;
parameter signed W59TO37 = 0;
parameter signed W59TO38 = 0;
parameter signed W59TO39 = 0;
parameter signed W59TO40 = 0;
parameter signed W59TO41 = 0;
parameter signed W59TO42 = 0;
parameter signed W59TO43 = 0;
parameter signed W59TO44 = 0;
parameter signed W59TO45 = 0;
parameter signed W59TO46 = 0;
parameter signed W59TO47 = 0;
parameter signed W59TO48 = 0;
parameter signed W59TO49 = 0;
parameter signed W59TO50 = 0;
parameter signed W59TO51 = 0;
parameter signed W59TO52 = 0;
parameter signed W59TO53 = 0;
parameter signed W59TO54 = 0;
parameter signed W59TO55 = 0;
parameter signed W59TO56 = 0;
parameter signed W59TO57 = 0;
parameter signed W59TO58 = 0;
parameter signed W59TO59 = 0;
parameter signed W59TO60 = 0;
parameter signed W59TO61 = 0;
parameter signed W59TO62 = 0;
parameter signed W59TO63 = 0;
parameter signed W60TO0 = 0;
parameter signed W60TO1 = 0;
parameter signed W60TO2 = 0;
parameter signed W60TO3 = 0;
parameter signed W60TO4 = 0;
parameter signed W60TO5 = 0;
parameter signed W60TO6 = 0;
parameter signed W60TO7 = 0;
parameter signed W60TO8 = 0;
parameter signed W60TO9 = 0;
parameter signed W60TO10 = 0;
parameter signed W60TO11 = 0;
parameter signed W60TO12 = 0;
parameter signed W60TO13 = 0;
parameter signed W60TO14 = 0;
parameter signed W60TO15 = 0;
parameter signed W60TO16 = 0;
parameter signed W60TO17 = 0;
parameter signed W60TO18 = 0;
parameter signed W60TO19 = 0;
parameter signed W60TO20 = 0;
parameter signed W60TO21 = 0;
parameter signed W60TO22 = 0;
parameter signed W60TO23 = 0;
parameter signed W60TO24 = 0;
parameter signed W60TO25 = 0;
parameter signed W60TO26 = 0;
parameter signed W60TO27 = 0;
parameter signed W60TO28 = 0;
parameter signed W60TO29 = 0;
parameter signed W60TO30 = 0;
parameter signed W60TO31 = 0;
parameter signed W60TO32 = 0;
parameter signed W60TO33 = 0;
parameter signed W60TO34 = 0;
parameter signed W60TO35 = 0;
parameter signed W60TO36 = 0;
parameter signed W60TO37 = 0;
parameter signed W60TO38 = 0;
parameter signed W60TO39 = 0;
parameter signed W60TO40 = 0;
parameter signed W60TO41 = 0;
parameter signed W60TO42 = 0;
parameter signed W60TO43 = 0;
parameter signed W60TO44 = 0;
parameter signed W60TO45 = 0;
parameter signed W60TO46 = 0;
parameter signed W60TO47 = 0;
parameter signed W60TO48 = 0;
parameter signed W60TO49 = 0;
parameter signed W60TO50 = 0;
parameter signed W60TO51 = 0;
parameter signed W60TO52 = 0;
parameter signed W60TO53 = 0;
parameter signed W60TO54 = 0;
parameter signed W60TO55 = 0;
parameter signed W60TO56 = 0;
parameter signed W60TO57 = 0;
parameter signed W60TO58 = 0;
parameter signed W60TO59 = 0;
parameter signed W60TO60 = 0;
parameter signed W60TO61 = 0;
parameter signed W60TO62 = 0;
parameter signed W60TO63 = 0;
parameter signed W61TO0 = 0;
parameter signed W61TO1 = 0;
parameter signed W61TO2 = 0;
parameter signed W61TO3 = 0;
parameter signed W61TO4 = 0;
parameter signed W61TO5 = 0;
parameter signed W61TO6 = 0;
parameter signed W61TO7 = 0;
parameter signed W61TO8 = 0;
parameter signed W61TO9 = 0;
parameter signed W61TO10 = 0;
parameter signed W61TO11 = 0;
parameter signed W61TO12 = 0;
parameter signed W61TO13 = 0;
parameter signed W61TO14 = 0;
parameter signed W61TO15 = 0;
parameter signed W61TO16 = 0;
parameter signed W61TO17 = 0;
parameter signed W61TO18 = 0;
parameter signed W61TO19 = 0;
parameter signed W61TO20 = 0;
parameter signed W61TO21 = 0;
parameter signed W61TO22 = 0;
parameter signed W61TO23 = 0;
parameter signed W61TO24 = 0;
parameter signed W61TO25 = 0;
parameter signed W61TO26 = 0;
parameter signed W61TO27 = 0;
parameter signed W61TO28 = 0;
parameter signed W61TO29 = 0;
parameter signed W61TO30 = 0;
parameter signed W61TO31 = 0;
parameter signed W61TO32 = 0;
parameter signed W61TO33 = 0;
parameter signed W61TO34 = 0;
parameter signed W61TO35 = 0;
parameter signed W61TO36 = 0;
parameter signed W61TO37 = 0;
parameter signed W61TO38 = 0;
parameter signed W61TO39 = 0;
parameter signed W61TO40 = 0;
parameter signed W61TO41 = 0;
parameter signed W61TO42 = 0;
parameter signed W61TO43 = 0;
parameter signed W61TO44 = 0;
parameter signed W61TO45 = 0;
parameter signed W61TO46 = 0;
parameter signed W61TO47 = 0;
parameter signed W61TO48 = 0;
parameter signed W61TO49 = 0;
parameter signed W61TO50 = 0;
parameter signed W61TO51 = 0;
parameter signed W61TO52 = 0;
parameter signed W61TO53 = 0;
parameter signed W61TO54 = 0;
parameter signed W61TO55 = 0;
parameter signed W61TO56 = 0;
parameter signed W61TO57 = 0;
parameter signed W61TO58 = 0;
parameter signed W61TO59 = 0;
parameter signed W61TO60 = 0;
parameter signed W61TO61 = 0;
parameter signed W61TO62 = 0;
parameter signed W61TO63 = 0;
parameter signed W62TO0 = 0;
parameter signed W62TO1 = 0;
parameter signed W62TO2 = 0;
parameter signed W62TO3 = 0;
parameter signed W62TO4 = 0;
parameter signed W62TO5 = 0;
parameter signed W62TO6 = 0;
parameter signed W62TO7 = 0;
parameter signed W62TO8 = 0;
parameter signed W62TO9 = 0;
parameter signed W62TO10 = 0;
parameter signed W62TO11 = 0;
parameter signed W62TO12 = 0;
parameter signed W62TO13 = 0;
parameter signed W62TO14 = 0;
parameter signed W62TO15 = 0;
parameter signed W62TO16 = 0;
parameter signed W62TO17 = 0;
parameter signed W62TO18 = 0;
parameter signed W62TO19 = 0;
parameter signed W62TO20 = 0;
parameter signed W62TO21 = 0;
parameter signed W62TO22 = 0;
parameter signed W62TO23 = 0;
parameter signed W62TO24 = 0;
parameter signed W62TO25 = 0;
parameter signed W62TO26 = 0;
parameter signed W62TO27 = 0;
parameter signed W62TO28 = 0;
parameter signed W62TO29 = 0;
parameter signed W62TO30 = 0;
parameter signed W62TO31 = 0;
parameter signed W62TO32 = 0;
parameter signed W62TO33 = 0;
parameter signed W62TO34 = 0;
parameter signed W62TO35 = 0;
parameter signed W62TO36 = 0;
parameter signed W62TO37 = 0;
parameter signed W62TO38 = 0;
parameter signed W62TO39 = 0;
parameter signed W62TO40 = 0;
parameter signed W62TO41 = 0;
parameter signed W62TO42 = 0;
parameter signed W62TO43 = 0;
parameter signed W62TO44 = 0;
parameter signed W62TO45 = 0;
parameter signed W62TO46 = 0;
parameter signed W62TO47 = 0;
parameter signed W62TO48 = 0;
parameter signed W62TO49 = 0;
parameter signed W62TO50 = 0;
parameter signed W62TO51 = 0;
parameter signed W62TO52 = 0;
parameter signed W62TO53 = 0;
parameter signed W62TO54 = 0;
parameter signed W62TO55 = 0;
parameter signed W62TO56 = 0;
parameter signed W62TO57 = 0;
parameter signed W62TO58 = 0;
parameter signed W62TO59 = 0;
parameter signed W62TO60 = 0;
parameter signed W62TO61 = 0;
parameter signed W62TO62 = 0;
parameter signed W62TO63 = 0;
parameter signed W63TO0 = 0;
parameter signed W63TO1 = 0;
parameter signed W63TO2 = 0;
parameter signed W63TO3 = 0;
parameter signed W63TO4 = 0;
parameter signed W63TO5 = 0;
parameter signed W63TO6 = 0;
parameter signed W63TO7 = 0;
parameter signed W63TO8 = 0;
parameter signed W63TO9 = 0;
parameter signed W63TO10 = 0;
parameter signed W63TO11 = 0;
parameter signed W63TO12 = 0;
parameter signed W63TO13 = 0;
parameter signed W63TO14 = 0;
parameter signed W63TO15 = 0;
parameter signed W63TO16 = 0;
parameter signed W63TO17 = 0;
parameter signed W63TO18 = 0;
parameter signed W63TO19 = 0;
parameter signed W63TO20 = 0;
parameter signed W63TO21 = 0;
parameter signed W63TO22 = 0;
parameter signed W63TO23 = 0;
parameter signed W63TO24 = 0;
parameter signed W63TO25 = 0;
parameter signed W63TO26 = 0;
parameter signed W63TO27 = 0;
parameter signed W63TO28 = 0;
parameter signed W63TO29 = 0;
parameter signed W63TO30 = 0;
parameter signed W63TO31 = 0;
parameter signed W63TO32 = 0;
parameter signed W63TO33 = 0;
parameter signed W63TO34 = 0;
parameter signed W63TO35 = 0;
parameter signed W63TO36 = 0;
parameter signed W63TO37 = 0;
parameter signed W63TO38 = 0;
parameter signed W63TO39 = 0;
parameter signed W63TO40 = 0;
parameter signed W63TO41 = 0;
parameter signed W63TO42 = 0;
parameter signed W63TO43 = 0;
parameter signed W63TO44 = 0;
parameter signed W63TO45 = 0;
parameter signed W63TO46 = 0;
parameter signed W63TO47 = 0;
parameter signed W63TO48 = 0;
parameter signed W63TO49 = 0;
parameter signed W63TO50 = 0;
parameter signed W63TO51 = 0;
parameter signed W63TO52 = 0;
parameter signed W63TO53 = 0;
parameter signed W63TO54 = 0;
parameter signed W63TO55 = 0;
parameter signed W63TO56 = 0;
parameter signed W63TO57 = 0;
parameter signed W63TO58 = 0;
parameter signed W63TO59 = 0;
parameter signed W63TO60 = 0;
parameter signed W63TO61 = 0;
parameter signed W63TO62 = 0;
parameter signed W63TO63 = 0;
parameter signed W64TO0 = 0;
parameter signed W64TO1 = 0;
parameter signed W64TO2 = 0;
parameter signed W64TO3 = 0;
parameter signed W64TO4 = 0;
parameter signed W64TO5 = 0;
parameter signed W64TO6 = 0;
parameter signed W64TO7 = 0;
parameter signed W64TO8 = 0;
parameter signed W64TO9 = 0;
parameter signed W64TO10 = 0;
parameter signed W64TO11 = 0;
parameter signed W64TO12 = 0;
parameter signed W64TO13 = 0;
parameter signed W64TO14 = 0;
parameter signed W64TO15 = 0;
parameter signed W64TO16 = 0;
parameter signed W64TO17 = 0;
parameter signed W64TO18 = 0;
parameter signed W64TO19 = 0;
parameter signed W64TO20 = 0;
parameter signed W64TO21 = 0;
parameter signed W64TO22 = 0;
parameter signed W64TO23 = 0;
parameter signed W64TO24 = 0;
parameter signed W64TO25 = 0;
parameter signed W64TO26 = 0;
parameter signed W64TO27 = 0;
parameter signed W64TO28 = 0;
parameter signed W64TO29 = 0;
parameter signed W64TO30 = 0;
parameter signed W64TO31 = 0;
parameter signed W64TO32 = 0;
parameter signed W64TO33 = 0;
parameter signed W64TO34 = 0;
parameter signed W64TO35 = 0;
parameter signed W64TO36 = 0;
parameter signed W64TO37 = 0;
parameter signed W64TO38 = 0;
parameter signed W64TO39 = 0;
parameter signed W64TO40 = 0;
parameter signed W64TO41 = 0;
parameter signed W64TO42 = 0;
parameter signed W64TO43 = 0;
parameter signed W64TO44 = 0;
parameter signed W64TO45 = 0;
parameter signed W64TO46 = 0;
parameter signed W64TO47 = 0;
parameter signed W64TO48 = 0;
parameter signed W64TO49 = 0;
parameter signed W64TO50 = 0;
parameter signed W64TO51 = 0;
parameter signed W64TO52 = 0;
parameter signed W64TO53 = 0;
parameter signed W64TO54 = 0;
parameter signed W64TO55 = 0;
parameter signed W64TO56 = 0;
parameter signed W64TO57 = 0;
parameter signed W64TO58 = 0;
parameter signed W64TO59 = 0;
parameter signed W64TO60 = 0;
parameter signed W64TO61 = 0;
parameter signed W64TO62 = 0;
parameter signed W64TO63 = 0;

input wire clk;
input wire rst;

input signed [15:0] in0;
input signed [15:0] in1;
input signed [15:0] in2;
input signed [15:0] in3;
input signed [15:0] in4;
input signed [15:0] in5;
input signed [15:0] in6;
input signed [15:0] in7;
input signed [15:0] in8;
input signed [15:0] in9;
input signed [15:0] in10;
input signed [15:0] in11;
input signed [15:0] in12;
input signed [15:0] in13;
input signed [15:0] in14;
input signed [15:0] in15;
input signed [15:0] in16;
input signed [15:0] in17;
input signed [15:0] in18;
input signed [15:0] in19;
input signed [15:0] in20;
input signed [15:0] in21;
input signed [15:0] in22;
input signed [15:0] in23;
input signed [15:0] in24;
input signed [15:0] in25;
input signed [15:0] in26;
input signed [15:0] in27;
input signed [15:0] in28;
input signed [15:0] in29;
input signed [15:0] in30;
input signed [15:0] in31;
input signed [15:0] in32;
input signed [15:0] in33;
input signed [15:0] in34;
input signed [15:0] in35;
input signed [15:0] in36;
input signed [15:0] in37;
input signed [15:0] in38;
input signed [15:0] in39;
input signed [15:0] in40;
input signed [15:0] in41;
input signed [15:0] in42;
input signed [15:0] in43;
input signed [15:0] in44;
input signed [15:0] in45;
input signed [15:0] in46;
input signed [15:0] in47;
input signed [15:0] in48;
input signed [15:0] in49;
input signed [15:0] in50;
input signed [15:0] in51;
input signed [15:0] in52;
input signed [15:0] in53;
input signed [15:0] in54;
input signed [15:0] in55;
input signed [15:0] in56;
input signed [15:0] in57;
input signed [15:0] in58;
input signed [15:0] in59;
input signed [15:0] in60;
input signed [15:0] in61;
input signed [15:0] in62;
input signed [15:0] in63;
input signed [15:0] in64;

output signed [15:0] out0;
output signed [15:0] out1;
output signed [15:0] out2;
output signed [15:0] out3;
output signed [15:0] out4;
output signed [15:0] out5;
output signed [15:0] out6;
output signed [15:0] out7;
output signed [15:0] out8;
output signed [15:0] out9;
output signed [15:0] out10;
output signed [15:0] out11;
output signed [15:0] out12;
output signed [15:0] out13;
output signed [15:0] out14;
output signed [15:0] out15;
output signed [15:0] out16;
output signed [15:0] out17;
output signed [15:0] out18;
output signed [15:0] out19;
output signed [15:0] out20;
output signed [15:0] out21;
output signed [15:0] out22;
output signed [15:0] out23;
output signed [15:0] out24;
output signed [15:0] out25;
output signed [15:0] out26;
output signed [15:0] out27;
output signed [15:0] out28;
output signed [15:0] out29;
output signed [15:0] out30;
output signed [15:0] out31;
output signed [15:0] out32;
output signed [15:0] out33;
output signed [15:0] out34;
output signed [15:0] out35;
output signed [15:0] out36;
output signed [15:0] out37;
output signed [15:0] out38;
output signed [15:0] out39;
output signed [15:0] out40;
output signed [15:0] out41;
output signed [15:0] out42;
output signed [15:0] out43;
output signed [15:0] out44;
output signed [15:0] out45;
output signed [15:0] out46;
output signed [15:0] out47;
output signed [15:0] out48;
output signed [15:0] out49;
output signed [15:0] out50;
output signed [15:0] out51;
output signed [15:0] out52;
output signed [15:0] out53;
output signed [15:0] out54;
output signed [15:0] out55;
output signed [15:0] out56;
output signed [15:0] out57;
output signed [15:0] out58;
output signed [15:0] out59;
output signed [15:0] out60;
output signed [15:0] out61;
output signed [15:0] out62;
output signed [15:0] out63;

neuron65in #(.BIAS(BIAS0), .W0(W0TO0), .W1(W1TO0), .W2(W2TO0), .W3(W3TO0), .W4(W4TO0), .W5(W5TO0), .W6(W6TO0), .W7(W7TO0), .W8(W8TO0), .W9(W9TO0), .W10(W10TO0), .W11(W11TO0), .W12(W12TO0), .W13(W13TO0), .W14(W14TO0), .W15(W15TO0), .W16(W16TO0), .W17(W17TO0), .W18(W18TO0), .W19(W19TO0), .W20(W20TO0), .W21(W21TO0), .W22(W22TO0), .W23(W23TO0), .W24(W24TO0), .W25(W25TO0), .W26(W26TO0), .W27(W27TO0), .W28(W28TO0), .W29(W29TO0), .W30(W30TO0), .W31(W31TO0), .W32(W32TO0), .W33(W33TO0), .W34(W34TO0), .W35(W35TO0), .W36(W36TO0), .W37(W37TO0), .W38(W38TO0), .W39(W39TO0), .W40(W40TO0), .W41(W41TO0), .W42(W42TO0), .W43(W43TO0), .W44(W44TO0), .W45(W45TO0), .W46(W46TO0), .W47(W47TO0), .W48(W48TO0), .W49(W49TO0), .W50(W50TO0), .W51(W51TO0), .W52(W52TO0), .W53(W53TO0), .W54(W54TO0), .W55(W55TO0), .W56(W56TO0), .W57(W57TO0), .W58(W58TO0), .W59(W59TO0), .W60(W60TO0), .W61(W61TO0), .W62(W62TO0), .W63(W63TO0), .W64(W64TO0)) neuron0(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out0));
neuron65in #(.BIAS(BIAS1), .W0(W0TO1), .W1(W1TO1), .W2(W2TO1), .W3(W3TO1), .W4(W4TO1), .W5(W5TO1), .W6(W6TO1), .W7(W7TO1), .W8(W8TO1), .W9(W9TO1), .W10(W10TO1), .W11(W11TO1), .W12(W12TO1), .W13(W13TO1), .W14(W14TO1), .W15(W15TO1), .W16(W16TO1), .W17(W17TO1), .W18(W18TO1), .W19(W19TO1), .W20(W20TO1), .W21(W21TO1), .W22(W22TO1), .W23(W23TO1), .W24(W24TO1), .W25(W25TO1), .W26(W26TO1), .W27(W27TO1), .W28(W28TO1), .W29(W29TO1), .W30(W30TO1), .W31(W31TO1), .W32(W32TO1), .W33(W33TO1), .W34(W34TO1), .W35(W35TO1), .W36(W36TO1), .W37(W37TO1), .W38(W38TO1), .W39(W39TO1), .W40(W40TO1), .W41(W41TO1), .W42(W42TO1), .W43(W43TO1), .W44(W44TO1), .W45(W45TO1), .W46(W46TO1), .W47(W47TO1), .W48(W48TO1), .W49(W49TO1), .W50(W50TO1), .W51(W51TO1), .W52(W52TO1), .W53(W53TO1), .W54(W54TO1), .W55(W55TO1), .W56(W56TO1), .W57(W57TO1), .W58(W58TO1), .W59(W59TO1), .W60(W60TO1), .W61(W61TO1), .W62(W62TO1), .W63(W63TO1), .W64(W64TO1)) neuron1(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out1));
neuron65in #(.BIAS(BIAS2), .W0(W0TO2), .W1(W1TO2), .W2(W2TO2), .W3(W3TO2), .W4(W4TO2), .W5(W5TO2), .W6(W6TO2), .W7(W7TO2), .W8(W8TO2), .W9(W9TO2), .W10(W10TO2), .W11(W11TO2), .W12(W12TO2), .W13(W13TO2), .W14(W14TO2), .W15(W15TO2), .W16(W16TO2), .W17(W17TO2), .W18(W18TO2), .W19(W19TO2), .W20(W20TO2), .W21(W21TO2), .W22(W22TO2), .W23(W23TO2), .W24(W24TO2), .W25(W25TO2), .W26(W26TO2), .W27(W27TO2), .W28(W28TO2), .W29(W29TO2), .W30(W30TO2), .W31(W31TO2), .W32(W32TO2), .W33(W33TO2), .W34(W34TO2), .W35(W35TO2), .W36(W36TO2), .W37(W37TO2), .W38(W38TO2), .W39(W39TO2), .W40(W40TO2), .W41(W41TO2), .W42(W42TO2), .W43(W43TO2), .W44(W44TO2), .W45(W45TO2), .W46(W46TO2), .W47(W47TO2), .W48(W48TO2), .W49(W49TO2), .W50(W50TO2), .W51(W51TO2), .W52(W52TO2), .W53(W53TO2), .W54(W54TO2), .W55(W55TO2), .W56(W56TO2), .W57(W57TO2), .W58(W58TO2), .W59(W59TO2), .W60(W60TO2), .W61(W61TO2), .W62(W62TO2), .W63(W63TO2), .W64(W64TO2)) neuron2(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out2));
neuron65in #(.BIAS(BIAS3), .W0(W0TO3), .W1(W1TO3), .W2(W2TO3), .W3(W3TO3), .W4(W4TO3), .W5(W5TO3), .W6(W6TO3), .W7(W7TO3), .W8(W8TO3), .W9(W9TO3), .W10(W10TO3), .W11(W11TO3), .W12(W12TO3), .W13(W13TO3), .W14(W14TO3), .W15(W15TO3), .W16(W16TO3), .W17(W17TO3), .W18(W18TO3), .W19(W19TO3), .W20(W20TO3), .W21(W21TO3), .W22(W22TO3), .W23(W23TO3), .W24(W24TO3), .W25(W25TO3), .W26(W26TO3), .W27(W27TO3), .W28(W28TO3), .W29(W29TO3), .W30(W30TO3), .W31(W31TO3), .W32(W32TO3), .W33(W33TO3), .W34(W34TO3), .W35(W35TO3), .W36(W36TO3), .W37(W37TO3), .W38(W38TO3), .W39(W39TO3), .W40(W40TO3), .W41(W41TO3), .W42(W42TO3), .W43(W43TO3), .W44(W44TO3), .W45(W45TO3), .W46(W46TO3), .W47(W47TO3), .W48(W48TO3), .W49(W49TO3), .W50(W50TO3), .W51(W51TO3), .W52(W52TO3), .W53(W53TO3), .W54(W54TO3), .W55(W55TO3), .W56(W56TO3), .W57(W57TO3), .W58(W58TO3), .W59(W59TO3), .W60(W60TO3), .W61(W61TO3), .W62(W62TO3), .W63(W63TO3), .W64(W64TO3)) neuron3(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out3));
neuron65in #(.BIAS(BIAS4), .W0(W0TO4), .W1(W1TO4), .W2(W2TO4), .W3(W3TO4), .W4(W4TO4), .W5(W5TO4), .W6(W6TO4), .W7(W7TO4), .W8(W8TO4), .W9(W9TO4), .W10(W10TO4), .W11(W11TO4), .W12(W12TO4), .W13(W13TO4), .W14(W14TO4), .W15(W15TO4), .W16(W16TO4), .W17(W17TO4), .W18(W18TO4), .W19(W19TO4), .W20(W20TO4), .W21(W21TO4), .W22(W22TO4), .W23(W23TO4), .W24(W24TO4), .W25(W25TO4), .W26(W26TO4), .W27(W27TO4), .W28(W28TO4), .W29(W29TO4), .W30(W30TO4), .W31(W31TO4), .W32(W32TO4), .W33(W33TO4), .W34(W34TO4), .W35(W35TO4), .W36(W36TO4), .W37(W37TO4), .W38(W38TO4), .W39(W39TO4), .W40(W40TO4), .W41(W41TO4), .W42(W42TO4), .W43(W43TO4), .W44(W44TO4), .W45(W45TO4), .W46(W46TO4), .W47(W47TO4), .W48(W48TO4), .W49(W49TO4), .W50(W50TO4), .W51(W51TO4), .W52(W52TO4), .W53(W53TO4), .W54(W54TO4), .W55(W55TO4), .W56(W56TO4), .W57(W57TO4), .W58(W58TO4), .W59(W59TO4), .W60(W60TO4), .W61(W61TO4), .W62(W62TO4), .W63(W63TO4), .W64(W64TO4)) neuron4(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out4));
neuron65in #(.BIAS(BIAS5), .W0(W0TO5), .W1(W1TO5), .W2(W2TO5), .W3(W3TO5), .W4(W4TO5), .W5(W5TO5), .W6(W6TO5), .W7(W7TO5), .W8(W8TO5), .W9(W9TO5), .W10(W10TO5), .W11(W11TO5), .W12(W12TO5), .W13(W13TO5), .W14(W14TO5), .W15(W15TO5), .W16(W16TO5), .W17(W17TO5), .W18(W18TO5), .W19(W19TO5), .W20(W20TO5), .W21(W21TO5), .W22(W22TO5), .W23(W23TO5), .W24(W24TO5), .W25(W25TO5), .W26(W26TO5), .W27(W27TO5), .W28(W28TO5), .W29(W29TO5), .W30(W30TO5), .W31(W31TO5), .W32(W32TO5), .W33(W33TO5), .W34(W34TO5), .W35(W35TO5), .W36(W36TO5), .W37(W37TO5), .W38(W38TO5), .W39(W39TO5), .W40(W40TO5), .W41(W41TO5), .W42(W42TO5), .W43(W43TO5), .W44(W44TO5), .W45(W45TO5), .W46(W46TO5), .W47(W47TO5), .W48(W48TO5), .W49(W49TO5), .W50(W50TO5), .W51(W51TO5), .W52(W52TO5), .W53(W53TO5), .W54(W54TO5), .W55(W55TO5), .W56(W56TO5), .W57(W57TO5), .W58(W58TO5), .W59(W59TO5), .W60(W60TO5), .W61(W61TO5), .W62(W62TO5), .W63(W63TO5), .W64(W64TO5)) neuron5(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out5));
neuron65in #(.BIAS(BIAS6), .W0(W0TO6), .W1(W1TO6), .W2(W2TO6), .W3(W3TO6), .W4(W4TO6), .W5(W5TO6), .W6(W6TO6), .W7(W7TO6), .W8(W8TO6), .W9(W9TO6), .W10(W10TO6), .W11(W11TO6), .W12(W12TO6), .W13(W13TO6), .W14(W14TO6), .W15(W15TO6), .W16(W16TO6), .W17(W17TO6), .W18(W18TO6), .W19(W19TO6), .W20(W20TO6), .W21(W21TO6), .W22(W22TO6), .W23(W23TO6), .W24(W24TO6), .W25(W25TO6), .W26(W26TO6), .W27(W27TO6), .W28(W28TO6), .W29(W29TO6), .W30(W30TO6), .W31(W31TO6), .W32(W32TO6), .W33(W33TO6), .W34(W34TO6), .W35(W35TO6), .W36(W36TO6), .W37(W37TO6), .W38(W38TO6), .W39(W39TO6), .W40(W40TO6), .W41(W41TO6), .W42(W42TO6), .W43(W43TO6), .W44(W44TO6), .W45(W45TO6), .W46(W46TO6), .W47(W47TO6), .W48(W48TO6), .W49(W49TO6), .W50(W50TO6), .W51(W51TO6), .W52(W52TO6), .W53(W53TO6), .W54(W54TO6), .W55(W55TO6), .W56(W56TO6), .W57(W57TO6), .W58(W58TO6), .W59(W59TO6), .W60(W60TO6), .W61(W61TO6), .W62(W62TO6), .W63(W63TO6), .W64(W64TO6)) neuron6(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out6));
neuron65in #(.BIAS(BIAS7), .W0(W0TO7), .W1(W1TO7), .W2(W2TO7), .W3(W3TO7), .W4(W4TO7), .W5(W5TO7), .W6(W6TO7), .W7(W7TO7), .W8(W8TO7), .W9(W9TO7), .W10(W10TO7), .W11(W11TO7), .W12(W12TO7), .W13(W13TO7), .W14(W14TO7), .W15(W15TO7), .W16(W16TO7), .W17(W17TO7), .W18(W18TO7), .W19(W19TO7), .W20(W20TO7), .W21(W21TO7), .W22(W22TO7), .W23(W23TO7), .W24(W24TO7), .W25(W25TO7), .W26(W26TO7), .W27(W27TO7), .W28(W28TO7), .W29(W29TO7), .W30(W30TO7), .W31(W31TO7), .W32(W32TO7), .W33(W33TO7), .W34(W34TO7), .W35(W35TO7), .W36(W36TO7), .W37(W37TO7), .W38(W38TO7), .W39(W39TO7), .W40(W40TO7), .W41(W41TO7), .W42(W42TO7), .W43(W43TO7), .W44(W44TO7), .W45(W45TO7), .W46(W46TO7), .W47(W47TO7), .W48(W48TO7), .W49(W49TO7), .W50(W50TO7), .W51(W51TO7), .W52(W52TO7), .W53(W53TO7), .W54(W54TO7), .W55(W55TO7), .W56(W56TO7), .W57(W57TO7), .W58(W58TO7), .W59(W59TO7), .W60(W60TO7), .W61(W61TO7), .W62(W62TO7), .W63(W63TO7), .W64(W64TO7)) neuron7(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out7));
neuron65in #(.BIAS(BIAS8), .W0(W0TO8), .W1(W1TO8), .W2(W2TO8), .W3(W3TO8), .W4(W4TO8), .W5(W5TO8), .W6(W6TO8), .W7(W7TO8), .W8(W8TO8), .W9(W9TO8), .W10(W10TO8), .W11(W11TO8), .W12(W12TO8), .W13(W13TO8), .W14(W14TO8), .W15(W15TO8), .W16(W16TO8), .W17(W17TO8), .W18(W18TO8), .W19(W19TO8), .W20(W20TO8), .W21(W21TO8), .W22(W22TO8), .W23(W23TO8), .W24(W24TO8), .W25(W25TO8), .W26(W26TO8), .W27(W27TO8), .W28(W28TO8), .W29(W29TO8), .W30(W30TO8), .W31(W31TO8), .W32(W32TO8), .W33(W33TO8), .W34(W34TO8), .W35(W35TO8), .W36(W36TO8), .W37(W37TO8), .W38(W38TO8), .W39(W39TO8), .W40(W40TO8), .W41(W41TO8), .W42(W42TO8), .W43(W43TO8), .W44(W44TO8), .W45(W45TO8), .W46(W46TO8), .W47(W47TO8), .W48(W48TO8), .W49(W49TO8), .W50(W50TO8), .W51(W51TO8), .W52(W52TO8), .W53(W53TO8), .W54(W54TO8), .W55(W55TO8), .W56(W56TO8), .W57(W57TO8), .W58(W58TO8), .W59(W59TO8), .W60(W60TO8), .W61(W61TO8), .W62(W62TO8), .W63(W63TO8), .W64(W64TO8)) neuron8(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out8));
neuron65in #(.BIAS(BIAS9), .W0(W0TO9), .W1(W1TO9), .W2(W2TO9), .W3(W3TO9), .W4(W4TO9), .W5(W5TO9), .W6(W6TO9), .W7(W7TO9), .W8(W8TO9), .W9(W9TO9), .W10(W10TO9), .W11(W11TO9), .W12(W12TO9), .W13(W13TO9), .W14(W14TO9), .W15(W15TO9), .W16(W16TO9), .W17(W17TO9), .W18(W18TO9), .W19(W19TO9), .W20(W20TO9), .W21(W21TO9), .W22(W22TO9), .W23(W23TO9), .W24(W24TO9), .W25(W25TO9), .W26(W26TO9), .W27(W27TO9), .W28(W28TO9), .W29(W29TO9), .W30(W30TO9), .W31(W31TO9), .W32(W32TO9), .W33(W33TO9), .W34(W34TO9), .W35(W35TO9), .W36(W36TO9), .W37(W37TO9), .W38(W38TO9), .W39(W39TO9), .W40(W40TO9), .W41(W41TO9), .W42(W42TO9), .W43(W43TO9), .W44(W44TO9), .W45(W45TO9), .W46(W46TO9), .W47(W47TO9), .W48(W48TO9), .W49(W49TO9), .W50(W50TO9), .W51(W51TO9), .W52(W52TO9), .W53(W53TO9), .W54(W54TO9), .W55(W55TO9), .W56(W56TO9), .W57(W57TO9), .W58(W58TO9), .W59(W59TO9), .W60(W60TO9), .W61(W61TO9), .W62(W62TO9), .W63(W63TO9), .W64(W64TO9)) neuron9(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out9));
neuron65in #(.BIAS(BIAS10), .W0(W0TO10), .W1(W1TO10), .W2(W2TO10), .W3(W3TO10), .W4(W4TO10), .W5(W5TO10), .W6(W6TO10), .W7(W7TO10), .W8(W8TO10), .W9(W9TO10), .W10(W10TO10), .W11(W11TO10), .W12(W12TO10), .W13(W13TO10), .W14(W14TO10), .W15(W15TO10), .W16(W16TO10), .W17(W17TO10), .W18(W18TO10), .W19(W19TO10), .W20(W20TO10), .W21(W21TO10), .W22(W22TO10), .W23(W23TO10), .W24(W24TO10), .W25(W25TO10), .W26(W26TO10), .W27(W27TO10), .W28(W28TO10), .W29(W29TO10), .W30(W30TO10), .W31(W31TO10), .W32(W32TO10), .W33(W33TO10), .W34(W34TO10), .W35(W35TO10), .W36(W36TO10), .W37(W37TO10), .W38(W38TO10), .W39(W39TO10), .W40(W40TO10), .W41(W41TO10), .W42(W42TO10), .W43(W43TO10), .W44(W44TO10), .W45(W45TO10), .W46(W46TO10), .W47(W47TO10), .W48(W48TO10), .W49(W49TO10), .W50(W50TO10), .W51(W51TO10), .W52(W52TO10), .W53(W53TO10), .W54(W54TO10), .W55(W55TO10), .W56(W56TO10), .W57(W57TO10), .W58(W58TO10), .W59(W59TO10), .W60(W60TO10), .W61(W61TO10), .W62(W62TO10), .W63(W63TO10), .W64(W64TO10)) neuron10(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out10));
neuron65in #(.BIAS(BIAS11), .W0(W0TO11), .W1(W1TO11), .W2(W2TO11), .W3(W3TO11), .W4(W4TO11), .W5(W5TO11), .W6(W6TO11), .W7(W7TO11), .W8(W8TO11), .W9(W9TO11), .W10(W10TO11), .W11(W11TO11), .W12(W12TO11), .W13(W13TO11), .W14(W14TO11), .W15(W15TO11), .W16(W16TO11), .W17(W17TO11), .W18(W18TO11), .W19(W19TO11), .W20(W20TO11), .W21(W21TO11), .W22(W22TO11), .W23(W23TO11), .W24(W24TO11), .W25(W25TO11), .W26(W26TO11), .W27(W27TO11), .W28(W28TO11), .W29(W29TO11), .W30(W30TO11), .W31(W31TO11), .W32(W32TO11), .W33(W33TO11), .W34(W34TO11), .W35(W35TO11), .W36(W36TO11), .W37(W37TO11), .W38(W38TO11), .W39(W39TO11), .W40(W40TO11), .W41(W41TO11), .W42(W42TO11), .W43(W43TO11), .W44(W44TO11), .W45(W45TO11), .W46(W46TO11), .W47(W47TO11), .W48(W48TO11), .W49(W49TO11), .W50(W50TO11), .W51(W51TO11), .W52(W52TO11), .W53(W53TO11), .W54(W54TO11), .W55(W55TO11), .W56(W56TO11), .W57(W57TO11), .W58(W58TO11), .W59(W59TO11), .W60(W60TO11), .W61(W61TO11), .W62(W62TO11), .W63(W63TO11), .W64(W64TO11)) neuron11(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out11));
neuron65in #(.BIAS(BIAS12), .W0(W0TO12), .W1(W1TO12), .W2(W2TO12), .W3(W3TO12), .W4(W4TO12), .W5(W5TO12), .W6(W6TO12), .W7(W7TO12), .W8(W8TO12), .W9(W9TO12), .W10(W10TO12), .W11(W11TO12), .W12(W12TO12), .W13(W13TO12), .W14(W14TO12), .W15(W15TO12), .W16(W16TO12), .W17(W17TO12), .W18(W18TO12), .W19(W19TO12), .W20(W20TO12), .W21(W21TO12), .W22(W22TO12), .W23(W23TO12), .W24(W24TO12), .W25(W25TO12), .W26(W26TO12), .W27(W27TO12), .W28(W28TO12), .W29(W29TO12), .W30(W30TO12), .W31(W31TO12), .W32(W32TO12), .W33(W33TO12), .W34(W34TO12), .W35(W35TO12), .W36(W36TO12), .W37(W37TO12), .W38(W38TO12), .W39(W39TO12), .W40(W40TO12), .W41(W41TO12), .W42(W42TO12), .W43(W43TO12), .W44(W44TO12), .W45(W45TO12), .W46(W46TO12), .W47(W47TO12), .W48(W48TO12), .W49(W49TO12), .W50(W50TO12), .W51(W51TO12), .W52(W52TO12), .W53(W53TO12), .W54(W54TO12), .W55(W55TO12), .W56(W56TO12), .W57(W57TO12), .W58(W58TO12), .W59(W59TO12), .W60(W60TO12), .W61(W61TO12), .W62(W62TO12), .W63(W63TO12), .W64(W64TO12)) neuron12(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out12));
neuron65in #(.BIAS(BIAS13), .W0(W0TO13), .W1(W1TO13), .W2(W2TO13), .W3(W3TO13), .W4(W4TO13), .W5(W5TO13), .W6(W6TO13), .W7(W7TO13), .W8(W8TO13), .W9(W9TO13), .W10(W10TO13), .W11(W11TO13), .W12(W12TO13), .W13(W13TO13), .W14(W14TO13), .W15(W15TO13), .W16(W16TO13), .W17(W17TO13), .W18(W18TO13), .W19(W19TO13), .W20(W20TO13), .W21(W21TO13), .W22(W22TO13), .W23(W23TO13), .W24(W24TO13), .W25(W25TO13), .W26(W26TO13), .W27(W27TO13), .W28(W28TO13), .W29(W29TO13), .W30(W30TO13), .W31(W31TO13), .W32(W32TO13), .W33(W33TO13), .W34(W34TO13), .W35(W35TO13), .W36(W36TO13), .W37(W37TO13), .W38(W38TO13), .W39(W39TO13), .W40(W40TO13), .W41(W41TO13), .W42(W42TO13), .W43(W43TO13), .W44(W44TO13), .W45(W45TO13), .W46(W46TO13), .W47(W47TO13), .W48(W48TO13), .W49(W49TO13), .W50(W50TO13), .W51(W51TO13), .W52(W52TO13), .W53(W53TO13), .W54(W54TO13), .W55(W55TO13), .W56(W56TO13), .W57(W57TO13), .W58(W58TO13), .W59(W59TO13), .W60(W60TO13), .W61(W61TO13), .W62(W62TO13), .W63(W63TO13), .W64(W64TO13)) neuron13(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out13));
neuron65in #(.BIAS(BIAS14), .W0(W0TO14), .W1(W1TO14), .W2(W2TO14), .W3(W3TO14), .W4(W4TO14), .W5(W5TO14), .W6(W6TO14), .W7(W7TO14), .W8(W8TO14), .W9(W9TO14), .W10(W10TO14), .W11(W11TO14), .W12(W12TO14), .W13(W13TO14), .W14(W14TO14), .W15(W15TO14), .W16(W16TO14), .W17(W17TO14), .W18(W18TO14), .W19(W19TO14), .W20(W20TO14), .W21(W21TO14), .W22(W22TO14), .W23(W23TO14), .W24(W24TO14), .W25(W25TO14), .W26(W26TO14), .W27(W27TO14), .W28(W28TO14), .W29(W29TO14), .W30(W30TO14), .W31(W31TO14), .W32(W32TO14), .W33(W33TO14), .W34(W34TO14), .W35(W35TO14), .W36(W36TO14), .W37(W37TO14), .W38(W38TO14), .W39(W39TO14), .W40(W40TO14), .W41(W41TO14), .W42(W42TO14), .W43(W43TO14), .W44(W44TO14), .W45(W45TO14), .W46(W46TO14), .W47(W47TO14), .W48(W48TO14), .W49(W49TO14), .W50(W50TO14), .W51(W51TO14), .W52(W52TO14), .W53(W53TO14), .W54(W54TO14), .W55(W55TO14), .W56(W56TO14), .W57(W57TO14), .W58(W58TO14), .W59(W59TO14), .W60(W60TO14), .W61(W61TO14), .W62(W62TO14), .W63(W63TO14), .W64(W64TO14)) neuron14(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out14));
neuron65in #(.BIAS(BIAS15), .W0(W0TO15), .W1(W1TO15), .W2(W2TO15), .W3(W3TO15), .W4(W4TO15), .W5(W5TO15), .W6(W6TO15), .W7(W7TO15), .W8(W8TO15), .W9(W9TO15), .W10(W10TO15), .W11(W11TO15), .W12(W12TO15), .W13(W13TO15), .W14(W14TO15), .W15(W15TO15), .W16(W16TO15), .W17(W17TO15), .W18(W18TO15), .W19(W19TO15), .W20(W20TO15), .W21(W21TO15), .W22(W22TO15), .W23(W23TO15), .W24(W24TO15), .W25(W25TO15), .W26(W26TO15), .W27(W27TO15), .W28(W28TO15), .W29(W29TO15), .W30(W30TO15), .W31(W31TO15), .W32(W32TO15), .W33(W33TO15), .W34(W34TO15), .W35(W35TO15), .W36(W36TO15), .W37(W37TO15), .W38(W38TO15), .W39(W39TO15), .W40(W40TO15), .W41(W41TO15), .W42(W42TO15), .W43(W43TO15), .W44(W44TO15), .W45(W45TO15), .W46(W46TO15), .W47(W47TO15), .W48(W48TO15), .W49(W49TO15), .W50(W50TO15), .W51(W51TO15), .W52(W52TO15), .W53(W53TO15), .W54(W54TO15), .W55(W55TO15), .W56(W56TO15), .W57(W57TO15), .W58(W58TO15), .W59(W59TO15), .W60(W60TO15), .W61(W61TO15), .W62(W62TO15), .W63(W63TO15), .W64(W64TO15)) neuron15(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out15));
neuron65in #(.BIAS(BIAS16), .W0(W0TO16), .W1(W1TO16), .W2(W2TO16), .W3(W3TO16), .W4(W4TO16), .W5(W5TO16), .W6(W6TO16), .W7(W7TO16), .W8(W8TO16), .W9(W9TO16), .W10(W10TO16), .W11(W11TO16), .W12(W12TO16), .W13(W13TO16), .W14(W14TO16), .W15(W15TO16), .W16(W16TO16), .W17(W17TO16), .W18(W18TO16), .W19(W19TO16), .W20(W20TO16), .W21(W21TO16), .W22(W22TO16), .W23(W23TO16), .W24(W24TO16), .W25(W25TO16), .W26(W26TO16), .W27(W27TO16), .W28(W28TO16), .W29(W29TO16), .W30(W30TO16), .W31(W31TO16), .W32(W32TO16), .W33(W33TO16), .W34(W34TO16), .W35(W35TO16), .W36(W36TO16), .W37(W37TO16), .W38(W38TO16), .W39(W39TO16), .W40(W40TO16), .W41(W41TO16), .W42(W42TO16), .W43(W43TO16), .W44(W44TO16), .W45(W45TO16), .W46(W46TO16), .W47(W47TO16), .W48(W48TO16), .W49(W49TO16), .W50(W50TO16), .W51(W51TO16), .W52(W52TO16), .W53(W53TO16), .W54(W54TO16), .W55(W55TO16), .W56(W56TO16), .W57(W57TO16), .W58(W58TO16), .W59(W59TO16), .W60(W60TO16), .W61(W61TO16), .W62(W62TO16), .W63(W63TO16), .W64(W64TO16)) neuron16(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out16));
neuron65in #(.BIAS(BIAS17), .W0(W0TO17), .W1(W1TO17), .W2(W2TO17), .W3(W3TO17), .W4(W4TO17), .W5(W5TO17), .W6(W6TO17), .W7(W7TO17), .W8(W8TO17), .W9(W9TO17), .W10(W10TO17), .W11(W11TO17), .W12(W12TO17), .W13(W13TO17), .W14(W14TO17), .W15(W15TO17), .W16(W16TO17), .W17(W17TO17), .W18(W18TO17), .W19(W19TO17), .W20(W20TO17), .W21(W21TO17), .W22(W22TO17), .W23(W23TO17), .W24(W24TO17), .W25(W25TO17), .W26(W26TO17), .W27(W27TO17), .W28(W28TO17), .W29(W29TO17), .W30(W30TO17), .W31(W31TO17), .W32(W32TO17), .W33(W33TO17), .W34(W34TO17), .W35(W35TO17), .W36(W36TO17), .W37(W37TO17), .W38(W38TO17), .W39(W39TO17), .W40(W40TO17), .W41(W41TO17), .W42(W42TO17), .W43(W43TO17), .W44(W44TO17), .W45(W45TO17), .W46(W46TO17), .W47(W47TO17), .W48(W48TO17), .W49(W49TO17), .W50(W50TO17), .W51(W51TO17), .W52(W52TO17), .W53(W53TO17), .W54(W54TO17), .W55(W55TO17), .W56(W56TO17), .W57(W57TO17), .W58(W58TO17), .W59(W59TO17), .W60(W60TO17), .W61(W61TO17), .W62(W62TO17), .W63(W63TO17), .W64(W64TO17)) neuron17(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out17));
neuron65in #(.BIAS(BIAS18), .W0(W0TO18), .W1(W1TO18), .W2(W2TO18), .W3(W3TO18), .W4(W4TO18), .W5(W5TO18), .W6(W6TO18), .W7(W7TO18), .W8(W8TO18), .W9(W9TO18), .W10(W10TO18), .W11(W11TO18), .W12(W12TO18), .W13(W13TO18), .W14(W14TO18), .W15(W15TO18), .W16(W16TO18), .W17(W17TO18), .W18(W18TO18), .W19(W19TO18), .W20(W20TO18), .W21(W21TO18), .W22(W22TO18), .W23(W23TO18), .W24(W24TO18), .W25(W25TO18), .W26(W26TO18), .W27(W27TO18), .W28(W28TO18), .W29(W29TO18), .W30(W30TO18), .W31(W31TO18), .W32(W32TO18), .W33(W33TO18), .W34(W34TO18), .W35(W35TO18), .W36(W36TO18), .W37(W37TO18), .W38(W38TO18), .W39(W39TO18), .W40(W40TO18), .W41(W41TO18), .W42(W42TO18), .W43(W43TO18), .W44(W44TO18), .W45(W45TO18), .W46(W46TO18), .W47(W47TO18), .W48(W48TO18), .W49(W49TO18), .W50(W50TO18), .W51(W51TO18), .W52(W52TO18), .W53(W53TO18), .W54(W54TO18), .W55(W55TO18), .W56(W56TO18), .W57(W57TO18), .W58(W58TO18), .W59(W59TO18), .W60(W60TO18), .W61(W61TO18), .W62(W62TO18), .W63(W63TO18), .W64(W64TO18)) neuron18(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out18));
neuron65in #(.BIAS(BIAS19), .W0(W0TO19), .W1(W1TO19), .W2(W2TO19), .W3(W3TO19), .W4(W4TO19), .W5(W5TO19), .W6(W6TO19), .W7(W7TO19), .W8(W8TO19), .W9(W9TO19), .W10(W10TO19), .W11(W11TO19), .W12(W12TO19), .W13(W13TO19), .W14(W14TO19), .W15(W15TO19), .W16(W16TO19), .W17(W17TO19), .W18(W18TO19), .W19(W19TO19), .W20(W20TO19), .W21(W21TO19), .W22(W22TO19), .W23(W23TO19), .W24(W24TO19), .W25(W25TO19), .W26(W26TO19), .W27(W27TO19), .W28(W28TO19), .W29(W29TO19), .W30(W30TO19), .W31(W31TO19), .W32(W32TO19), .W33(W33TO19), .W34(W34TO19), .W35(W35TO19), .W36(W36TO19), .W37(W37TO19), .W38(W38TO19), .W39(W39TO19), .W40(W40TO19), .W41(W41TO19), .W42(W42TO19), .W43(W43TO19), .W44(W44TO19), .W45(W45TO19), .W46(W46TO19), .W47(W47TO19), .W48(W48TO19), .W49(W49TO19), .W50(W50TO19), .W51(W51TO19), .W52(W52TO19), .W53(W53TO19), .W54(W54TO19), .W55(W55TO19), .W56(W56TO19), .W57(W57TO19), .W58(W58TO19), .W59(W59TO19), .W60(W60TO19), .W61(W61TO19), .W62(W62TO19), .W63(W63TO19), .W64(W64TO19)) neuron19(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out19));
neuron65in #(.BIAS(BIAS20), .W0(W0TO20), .W1(W1TO20), .W2(W2TO20), .W3(W3TO20), .W4(W4TO20), .W5(W5TO20), .W6(W6TO20), .W7(W7TO20), .W8(W8TO20), .W9(W9TO20), .W10(W10TO20), .W11(W11TO20), .W12(W12TO20), .W13(W13TO20), .W14(W14TO20), .W15(W15TO20), .W16(W16TO20), .W17(W17TO20), .W18(W18TO20), .W19(W19TO20), .W20(W20TO20), .W21(W21TO20), .W22(W22TO20), .W23(W23TO20), .W24(W24TO20), .W25(W25TO20), .W26(W26TO20), .W27(W27TO20), .W28(W28TO20), .W29(W29TO20), .W30(W30TO20), .W31(W31TO20), .W32(W32TO20), .W33(W33TO20), .W34(W34TO20), .W35(W35TO20), .W36(W36TO20), .W37(W37TO20), .W38(W38TO20), .W39(W39TO20), .W40(W40TO20), .W41(W41TO20), .W42(W42TO20), .W43(W43TO20), .W44(W44TO20), .W45(W45TO20), .W46(W46TO20), .W47(W47TO20), .W48(W48TO20), .W49(W49TO20), .W50(W50TO20), .W51(W51TO20), .W52(W52TO20), .W53(W53TO20), .W54(W54TO20), .W55(W55TO20), .W56(W56TO20), .W57(W57TO20), .W58(W58TO20), .W59(W59TO20), .W60(W60TO20), .W61(W61TO20), .W62(W62TO20), .W63(W63TO20), .W64(W64TO20)) neuron20(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out20));
neuron65in #(.BIAS(BIAS21), .W0(W0TO21), .W1(W1TO21), .W2(W2TO21), .W3(W3TO21), .W4(W4TO21), .W5(W5TO21), .W6(W6TO21), .W7(W7TO21), .W8(W8TO21), .W9(W9TO21), .W10(W10TO21), .W11(W11TO21), .W12(W12TO21), .W13(W13TO21), .W14(W14TO21), .W15(W15TO21), .W16(W16TO21), .W17(W17TO21), .W18(W18TO21), .W19(W19TO21), .W20(W20TO21), .W21(W21TO21), .W22(W22TO21), .W23(W23TO21), .W24(W24TO21), .W25(W25TO21), .W26(W26TO21), .W27(W27TO21), .W28(W28TO21), .W29(W29TO21), .W30(W30TO21), .W31(W31TO21), .W32(W32TO21), .W33(W33TO21), .W34(W34TO21), .W35(W35TO21), .W36(W36TO21), .W37(W37TO21), .W38(W38TO21), .W39(W39TO21), .W40(W40TO21), .W41(W41TO21), .W42(W42TO21), .W43(W43TO21), .W44(W44TO21), .W45(W45TO21), .W46(W46TO21), .W47(W47TO21), .W48(W48TO21), .W49(W49TO21), .W50(W50TO21), .W51(W51TO21), .W52(W52TO21), .W53(W53TO21), .W54(W54TO21), .W55(W55TO21), .W56(W56TO21), .W57(W57TO21), .W58(W58TO21), .W59(W59TO21), .W60(W60TO21), .W61(W61TO21), .W62(W62TO21), .W63(W63TO21), .W64(W64TO21)) neuron21(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out21));
neuron65in #(.BIAS(BIAS22), .W0(W0TO22), .W1(W1TO22), .W2(W2TO22), .W3(W3TO22), .W4(W4TO22), .W5(W5TO22), .W6(W6TO22), .W7(W7TO22), .W8(W8TO22), .W9(W9TO22), .W10(W10TO22), .W11(W11TO22), .W12(W12TO22), .W13(W13TO22), .W14(W14TO22), .W15(W15TO22), .W16(W16TO22), .W17(W17TO22), .W18(W18TO22), .W19(W19TO22), .W20(W20TO22), .W21(W21TO22), .W22(W22TO22), .W23(W23TO22), .W24(W24TO22), .W25(W25TO22), .W26(W26TO22), .W27(W27TO22), .W28(W28TO22), .W29(W29TO22), .W30(W30TO22), .W31(W31TO22), .W32(W32TO22), .W33(W33TO22), .W34(W34TO22), .W35(W35TO22), .W36(W36TO22), .W37(W37TO22), .W38(W38TO22), .W39(W39TO22), .W40(W40TO22), .W41(W41TO22), .W42(W42TO22), .W43(W43TO22), .W44(W44TO22), .W45(W45TO22), .W46(W46TO22), .W47(W47TO22), .W48(W48TO22), .W49(W49TO22), .W50(W50TO22), .W51(W51TO22), .W52(W52TO22), .W53(W53TO22), .W54(W54TO22), .W55(W55TO22), .W56(W56TO22), .W57(W57TO22), .W58(W58TO22), .W59(W59TO22), .W60(W60TO22), .W61(W61TO22), .W62(W62TO22), .W63(W63TO22), .W64(W64TO22)) neuron22(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out22));
neuron65in #(.BIAS(BIAS23), .W0(W0TO23), .W1(W1TO23), .W2(W2TO23), .W3(W3TO23), .W4(W4TO23), .W5(W5TO23), .W6(W6TO23), .W7(W7TO23), .W8(W8TO23), .W9(W9TO23), .W10(W10TO23), .W11(W11TO23), .W12(W12TO23), .W13(W13TO23), .W14(W14TO23), .W15(W15TO23), .W16(W16TO23), .W17(W17TO23), .W18(W18TO23), .W19(W19TO23), .W20(W20TO23), .W21(W21TO23), .W22(W22TO23), .W23(W23TO23), .W24(W24TO23), .W25(W25TO23), .W26(W26TO23), .W27(W27TO23), .W28(W28TO23), .W29(W29TO23), .W30(W30TO23), .W31(W31TO23), .W32(W32TO23), .W33(W33TO23), .W34(W34TO23), .W35(W35TO23), .W36(W36TO23), .W37(W37TO23), .W38(W38TO23), .W39(W39TO23), .W40(W40TO23), .W41(W41TO23), .W42(W42TO23), .W43(W43TO23), .W44(W44TO23), .W45(W45TO23), .W46(W46TO23), .W47(W47TO23), .W48(W48TO23), .W49(W49TO23), .W50(W50TO23), .W51(W51TO23), .W52(W52TO23), .W53(W53TO23), .W54(W54TO23), .W55(W55TO23), .W56(W56TO23), .W57(W57TO23), .W58(W58TO23), .W59(W59TO23), .W60(W60TO23), .W61(W61TO23), .W62(W62TO23), .W63(W63TO23), .W64(W64TO23)) neuron23(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out23));
neuron65in #(.BIAS(BIAS24), .W0(W0TO24), .W1(W1TO24), .W2(W2TO24), .W3(W3TO24), .W4(W4TO24), .W5(W5TO24), .W6(W6TO24), .W7(W7TO24), .W8(W8TO24), .W9(W9TO24), .W10(W10TO24), .W11(W11TO24), .W12(W12TO24), .W13(W13TO24), .W14(W14TO24), .W15(W15TO24), .W16(W16TO24), .W17(W17TO24), .W18(W18TO24), .W19(W19TO24), .W20(W20TO24), .W21(W21TO24), .W22(W22TO24), .W23(W23TO24), .W24(W24TO24), .W25(W25TO24), .W26(W26TO24), .W27(W27TO24), .W28(W28TO24), .W29(W29TO24), .W30(W30TO24), .W31(W31TO24), .W32(W32TO24), .W33(W33TO24), .W34(W34TO24), .W35(W35TO24), .W36(W36TO24), .W37(W37TO24), .W38(W38TO24), .W39(W39TO24), .W40(W40TO24), .W41(W41TO24), .W42(W42TO24), .W43(W43TO24), .W44(W44TO24), .W45(W45TO24), .W46(W46TO24), .W47(W47TO24), .W48(W48TO24), .W49(W49TO24), .W50(W50TO24), .W51(W51TO24), .W52(W52TO24), .W53(W53TO24), .W54(W54TO24), .W55(W55TO24), .W56(W56TO24), .W57(W57TO24), .W58(W58TO24), .W59(W59TO24), .W60(W60TO24), .W61(W61TO24), .W62(W62TO24), .W63(W63TO24), .W64(W64TO24)) neuron24(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out24));
neuron65in #(.BIAS(BIAS25), .W0(W0TO25), .W1(W1TO25), .W2(W2TO25), .W3(W3TO25), .W4(W4TO25), .W5(W5TO25), .W6(W6TO25), .W7(W7TO25), .W8(W8TO25), .W9(W9TO25), .W10(W10TO25), .W11(W11TO25), .W12(W12TO25), .W13(W13TO25), .W14(W14TO25), .W15(W15TO25), .W16(W16TO25), .W17(W17TO25), .W18(W18TO25), .W19(W19TO25), .W20(W20TO25), .W21(W21TO25), .W22(W22TO25), .W23(W23TO25), .W24(W24TO25), .W25(W25TO25), .W26(W26TO25), .W27(W27TO25), .W28(W28TO25), .W29(W29TO25), .W30(W30TO25), .W31(W31TO25), .W32(W32TO25), .W33(W33TO25), .W34(W34TO25), .W35(W35TO25), .W36(W36TO25), .W37(W37TO25), .W38(W38TO25), .W39(W39TO25), .W40(W40TO25), .W41(W41TO25), .W42(W42TO25), .W43(W43TO25), .W44(W44TO25), .W45(W45TO25), .W46(W46TO25), .W47(W47TO25), .W48(W48TO25), .W49(W49TO25), .W50(W50TO25), .W51(W51TO25), .W52(W52TO25), .W53(W53TO25), .W54(W54TO25), .W55(W55TO25), .W56(W56TO25), .W57(W57TO25), .W58(W58TO25), .W59(W59TO25), .W60(W60TO25), .W61(W61TO25), .W62(W62TO25), .W63(W63TO25), .W64(W64TO25)) neuron25(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out25));
neuron65in #(.BIAS(BIAS26), .W0(W0TO26), .W1(W1TO26), .W2(W2TO26), .W3(W3TO26), .W4(W4TO26), .W5(W5TO26), .W6(W6TO26), .W7(W7TO26), .W8(W8TO26), .W9(W9TO26), .W10(W10TO26), .W11(W11TO26), .W12(W12TO26), .W13(W13TO26), .W14(W14TO26), .W15(W15TO26), .W16(W16TO26), .W17(W17TO26), .W18(W18TO26), .W19(W19TO26), .W20(W20TO26), .W21(W21TO26), .W22(W22TO26), .W23(W23TO26), .W24(W24TO26), .W25(W25TO26), .W26(W26TO26), .W27(W27TO26), .W28(W28TO26), .W29(W29TO26), .W30(W30TO26), .W31(W31TO26), .W32(W32TO26), .W33(W33TO26), .W34(W34TO26), .W35(W35TO26), .W36(W36TO26), .W37(W37TO26), .W38(W38TO26), .W39(W39TO26), .W40(W40TO26), .W41(W41TO26), .W42(W42TO26), .W43(W43TO26), .W44(W44TO26), .W45(W45TO26), .W46(W46TO26), .W47(W47TO26), .W48(W48TO26), .W49(W49TO26), .W50(W50TO26), .W51(W51TO26), .W52(W52TO26), .W53(W53TO26), .W54(W54TO26), .W55(W55TO26), .W56(W56TO26), .W57(W57TO26), .W58(W58TO26), .W59(W59TO26), .W60(W60TO26), .W61(W61TO26), .W62(W62TO26), .W63(W63TO26), .W64(W64TO26)) neuron26(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out26));
neuron65in #(.BIAS(BIAS27), .W0(W0TO27), .W1(W1TO27), .W2(W2TO27), .W3(W3TO27), .W4(W4TO27), .W5(W5TO27), .W6(W6TO27), .W7(W7TO27), .W8(W8TO27), .W9(W9TO27), .W10(W10TO27), .W11(W11TO27), .W12(W12TO27), .W13(W13TO27), .W14(W14TO27), .W15(W15TO27), .W16(W16TO27), .W17(W17TO27), .W18(W18TO27), .W19(W19TO27), .W20(W20TO27), .W21(W21TO27), .W22(W22TO27), .W23(W23TO27), .W24(W24TO27), .W25(W25TO27), .W26(W26TO27), .W27(W27TO27), .W28(W28TO27), .W29(W29TO27), .W30(W30TO27), .W31(W31TO27), .W32(W32TO27), .W33(W33TO27), .W34(W34TO27), .W35(W35TO27), .W36(W36TO27), .W37(W37TO27), .W38(W38TO27), .W39(W39TO27), .W40(W40TO27), .W41(W41TO27), .W42(W42TO27), .W43(W43TO27), .W44(W44TO27), .W45(W45TO27), .W46(W46TO27), .W47(W47TO27), .W48(W48TO27), .W49(W49TO27), .W50(W50TO27), .W51(W51TO27), .W52(W52TO27), .W53(W53TO27), .W54(W54TO27), .W55(W55TO27), .W56(W56TO27), .W57(W57TO27), .W58(W58TO27), .W59(W59TO27), .W60(W60TO27), .W61(W61TO27), .W62(W62TO27), .W63(W63TO27), .W64(W64TO27)) neuron27(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out27));
neuron65in #(.BIAS(BIAS28), .W0(W0TO28), .W1(W1TO28), .W2(W2TO28), .W3(W3TO28), .W4(W4TO28), .W5(W5TO28), .W6(W6TO28), .W7(W7TO28), .W8(W8TO28), .W9(W9TO28), .W10(W10TO28), .W11(W11TO28), .W12(W12TO28), .W13(W13TO28), .W14(W14TO28), .W15(W15TO28), .W16(W16TO28), .W17(W17TO28), .W18(W18TO28), .W19(W19TO28), .W20(W20TO28), .W21(W21TO28), .W22(W22TO28), .W23(W23TO28), .W24(W24TO28), .W25(W25TO28), .W26(W26TO28), .W27(W27TO28), .W28(W28TO28), .W29(W29TO28), .W30(W30TO28), .W31(W31TO28), .W32(W32TO28), .W33(W33TO28), .W34(W34TO28), .W35(W35TO28), .W36(W36TO28), .W37(W37TO28), .W38(W38TO28), .W39(W39TO28), .W40(W40TO28), .W41(W41TO28), .W42(W42TO28), .W43(W43TO28), .W44(W44TO28), .W45(W45TO28), .W46(W46TO28), .W47(W47TO28), .W48(W48TO28), .W49(W49TO28), .W50(W50TO28), .W51(W51TO28), .W52(W52TO28), .W53(W53TO28), .W54(W54TO28), .W55(W55TO28), .W56(W56TO28), .W57(W57TO28), .W58(W58TO28), .W59(W59TO28), .W60(W60TO28), .W61(W61TO28), .W62(W62TO28), .W63(W63TO28), .W64(W64TO28)) neuron28(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out28));
neuron65in #(.BIAS(BIAS29), .W0(W0TO29), .W1(W1TO29), .W2(W2TO29), .W3(W3TO29), .W4(W4TO29), .W5(W5TO29), .W6(W6TO29), .W7(W7TO29), .W8(W8TO29), .W9(W9TO29), .W10(W10TO29), .W11(W11TO29), .W12(W12TO29), .W13(W13TO29), .W14(W14TO29), .W15(W15TO29), .W16(W16TO29), .W17(W17TO29), .W18(W18TO29), .W19(W19TO29), .W20(W20TO29), .W21(W21TO29), .W22(W22TO29), .W23(W23TO29), .W24(W24TO29), .W25(W25TO29), .W26(W26TO29), .W27(W27TO29), .W28(W28TO29), .W29(W29TO29), .W30(W30TO29), .W31(W31TO29), .W32(W32TO29), .W33(W33TO29), .W34(W34TO29), .W35(W35TO29), .W36(W36TO29), .W37(W37TO29), .W38(W38TO29), .W39(W39TO29), .W40(W40TO29), .W41(W41TO29), .W42(W42TO29), .W43(W43TO29), .W44(W44TO29), .W45(W45TO29), .W46(W46TO29), .W47(W47TO29), .W48(W48TO29), .W49(W49TO29), .W50(W50TO29), .W51(W51TO29), .W52(W52TO29), .W53(W53TO29), .W54(W54TO29), .W55(W55TO29), .W56(W56TO29), .W57(W57TO29), .W58(W58TO29), .W59(W59TO29), .W60(W60TO29), .W61(W61TO29), .W62(W62TO29), .W63(W63TO29), .W64(W64TO29)) neuron29(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out29));
neuron65in #(.BIAS(BIAS30), .W0(W0TO30), .W1(W1TO30), .W2(W2TO30), .W3(W3TO30), .W4(W4TO30), .W5(W5TO30), .W6(W6TO30), .W7(W7TO30), .W8(W8TO30), .W9(W9TO30), .W10(W10TO30), .W11(W11TO30), .W12(W12TO30), .W13(W13TO30), .W14(W14TO30), .W15(W15TO30), .W16(W16TO30), .W17(W17TO30), .W18(W18TO30), .W19(W19TO30), .W20(W20TO30), .W21(W21TO30), .W22(W22TO30), .W23(W23TO30), .W24(W24TO30), .W25(W25TO30), .W26(W26TO30), .W27(W27TO30), .W28(W28TO30), .W29(W29TO30), .W30(W30TO30), .W31(W31TO30), .W32(W32TO30), .W33(W33TO30), .W34(W34TO30), .W35(W35TO30), .W36(W36TO30), .W37(W37TO30), .W38(W38TO30), .W39(W39TO30), .W40(W40TO30), .W41(W41TO30), .W42(W42TO30), .W43(W43TO30), .W44(W44TO30), .W45(W45TO30), .W46(W46TO30), .W47(W47TO30), .W48(W48TO30), .W49(W49TO30), .W50(W50TO30), .W51(W51TO30), .W52(W52TO30), .W53(W53TO30), .W54(W54TO30), .W55(W55TO30), .W56(W56TO30), .W57(W57TO30), .W58(W58TO30), .W59(W59TO30), .W60(W60TO30), .W61(W61TO30), .W62(W62TO30), .W63(W63TO30), .W64(W64TO30)) neuron30(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out30));
neuron65in #(.BIAS(BIAS31), .W0(W0TO31), .W1(W1TO31), .W2(W2TO31), .W3(W3TO31), .W4(W4TO31), .W5(W5TO31), .W6(W6TO31), .W7(W7TO31), .W8(W8TO31), .W9(W9TO31), .W10(W10TO31), .W11(W11TO31), .W12(W12TO31), .W13(W13TO31), .W14(W14TO31), .W15(W15TO31), .W16(W16TO31), .W17(W17TO31), .W18(W18TO31), .W19(W19TO31), .W20(W20TO31), .W21(W21TO31), .W22(W22TO31), .W23(W23TO31), .W24(W24TO31), .W25(W25TO31), .W26(W26TO31), .W27(W27TO31), .W28(W28TO31), .W29(W29TO31), .W30(W30TO31), .W31(W31TO31), .W32(W32TO31), .W33(W33TO31), .W34(W34TO31), .W35(W35TO31), .W36(W36TO31), .W37(W37TO31), .W38(W38TO31), .W39(W39TO31), .W40(W40TO31), .W41(W41TO31), .W42(W42TO31), .W43(W43TO31), .W44(W44TO31), .W45(W45TO31), .W46(W46TO31), .W47(W47TO31), .W48(W48TO31), .W49(W49TO31), .W50(W50TO31), .W51(W51TO31), .W52(W52TO31), .W53(W53TO31), .W54(W54TO31), .W55(W55TO31), .W56(W56TO31), .W57(W57TO31), .W58(W58TO31), .W59(W59TO31), .W60(W60TO31), .W61(W61TO31), .W62(W62TO31), .W63(W63TO31), .W64(W64TO31)) neuron31(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out31));
neuron65in #(.BIAS(BIAS32), .W0(W0TO32), .W1(W1TO32), .W2(W2TO32), .W3(W3TO32), .W4(W4TO32), .W5(W5TO32), .W6(W6TO32), .W7(W7TO32), .W8(W8TO32), .W9(W9TO32), .W10(W10TO32), .W11(W11TO32), .W12(W12TO32), .W13(W13TO32), .W14(W14TO32), .W15(W15TO32), .W16(W16TO32), .W17(W17TO32), .W18(W18TO32), .W19(W19TO32), .W20(W20TO32), .W21(W21TO32), .W22(W22TO32), .W23(W23TO32), .W24(W24TO32), .W25(W25TO32), .W26(W26TO32), .W27(W27TO32), .W28(W28TO32), .W29(W29TO32), .W30(W30TO32), .W31(W31TO32), .W32(W32TO32), .W33(W33TO32), .W34(W34TO32), .W35(W35TO32), .W36(W36TO32), .W37(W37TO32), .W38(W38TO32), .W39(W39TO32), .W40(W40TO32), .W41(W41TO32), .W42(W42TO32), .W43(W43TO32), .W44(W44TO32), .W45(W45TO32), .W46(W46TO32), .W47(W47TO32), .W48(W48TO32), .W49(W49TO32), .W50(W50TO32), .W51(W51TO32), .W52(W52TO32), .W53(W53TO32), .W54(W54TO32), .W55(W55TO32), .W56(W56TO32), .W57(W57TO32), .W58(W58TO32), .W59(W59TO32), .W60(W60TO32), .W61(W61TO32), .W62(W62TO32), .W63(W63TO32), .W64(W64TO32)) neuron32(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out32));
neuron65in #(.BIAS(BIAS33), .W0(W0TO33), .W1(W1TO33), .W2(W2TO33), .W3(W3TO33), .W4(W4TO33), .W5(W5TO33), .W6(W6TO33), .W7(W7TO33), .W8(W8TO33), .W9(W9TO33), .W10(W10TO33), .W11(W11TO33), .W12(W12TO33), .W13(W13TO33), .W14(W14TO33), .W15(W15TO33), .W16(W16TO33), .W17(W17TO33), .W18(W18TO33), .W19(W19TO33), .W20(W20TO33), .W21(W21TO33), .W22(W22TO33), .W23(W23TO33), .W24(W24TO33), .W25(W25TO33), .W26(W26TO33), .W27(W27TO33), .W28(W28TO33), .W29(W29TO33), .W30(W30TO33), .W31(W31TO33), .W32(W32TO33), .W33(W33TO33), .W34(W34TO33), .W35(W35TO33), .W36(W36TO33), .W37(W37TO33), .W38(W38TO33), .W39(W39TO33), .W40(W40TO33), .W41(W41TO33), .W42(W42TO33), .W43(W43TO33), .W44(W44TO33), .W45(W45TO33), .W46(W46TO33), .W47(W47TO33), .W48(W48TO33), .W49(W49TO33), .W50(W50TO33), .W51(W51TO33), .W52(W52TO33), .W53(W53TO33), .W54(W54TO33), .W55(W55TO33), .W56(W56TO33), .W57(W57TO33), .W58(W58TO33), .W59(W59TO33), .W60(W60TO33), .W61(W61TO33), .W62(W62TO33), .W63(W63TO33), .W64(W64TO33)) neuron33(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out33));
neuron65in #(.BIAS(BIAS34), .W0(W0TO34), .W1(W1TO34), .W2(W2TO34), .W3(W3TO34), .W4(W4TO34), .W5(W5TO34), .W6(W6TO34), .W7(W7TO34), .W8(W8TO34), .W9(W9TO34), .W10(W10TO34), .W11(W11TO34), .W12(W12TO34), .W13(W13TO34), .W14(W14TO34), .W15(W15TO34), .W16(W16TO34), .W17(W17TO34), .W18(W18TO34), .W19(W19TO34), .W20(W20TO34), .W21(W21TO34), .W22(W22TO34), .W23(W23TO34), .W24(W24TO34), .W25(W25TO34), .W26(W26TO34), .W27(W27TO34), .W28(W28TO34), .W29(W29TO34), .W30(W30TO34), .W31(W31TO34), .W32(W32TO34), .W33(W33TO34), .W34(W34TO34), .W35(W35TO34), .W36(W36TO34), .W37(W37TO34), .W38(W38TO34), .W39(W39TO34), .W40(W40TO34), .W41(W41TO34), .W42(W42TO34), .W43(W43TO34), .W44(W44TO34), .W45(W45TO34), .W46(W46TO34), .W47(W47TO34), .W48(W48TO34), .W49(W49TO34), .W50(W50TO34), .W51(W51TO34), .W52(W52TO34), .W53(W53TO34), .W54(W54TO34), .W55(W55TO34), .W56(W56TO34), .W57(W57TO34), .W58(W58TO34), .W59(W59TO34), .W60(W60TO34), .W61(W61TO34), .W62(W62TO34), .W63(W63TO34), .W64(W64TO34)) neuron34(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out34));
neuron65in #(.BIAS(BIAS35), .W0(W0TO35), .W1(W1TO35), .W2(W2TO35), .W3(W3TO35), .W4(W4TO35), .W5(W5TO35), .W6(W6TO35), .W7(W7TO35), .W8(W8TO35), .W9(W9TO35), .W10(W10TO35), .W11(W11TO35), .W12(W12TO35), .W13(W13TO35), .W14(W14TO35), .W15(W15TO35), .W16(W16TO35), .W17(W17TO35), .W18(W18TO35), .W19(W19TO35), .W20(W20TO35), .W21(W21TO35), .W22(W22TO35), .W23(W23TO35), .W24(W24TO35), .W25(W25TO35), .W26(W26TO35), .W27(W27TO35), .W28(W28TO35), .W29(W29TO35), .W30(W30TO35), .W31(W31TO35), .W32(W32TO35), .W33(W33TO35), .W34(W34TO35), .W35(W35TO35), .W36(W36TO35), .W37(W37TO35), .W38(W38TO35), .W39(W39TO35), .W40(W40TO35), .W41(W41TO35), .W42(W42TO35), .W43(W43TO35), .W44(W44TO35), .W45(W45TO35), .W46(W46TO35), .W47(W47TO35), .W48(W48TO35), .W49(W49TO35), .W50(W50TO35), .W51(W51TO35), .W52(W52TO35), .W53(W53TO35), .W54(W54TO35), .W55(W55TO35), .W56(W56TO35), .W57(W57TO35), .W58(W58TO35), .W59(W59TO35), .W60(W60TO35), .W61(W61TO35), .W62(W62TO35), .W63(W63TO35), .W64(W64TO35)) neuron35(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out35));
neuron65in #(.BIAS(BIAS36), .W0(W0TO36), .W1(W1TO36), .W2(W2TO36), .W3(W3TO36), .W4(W4TO36), .W5(W5TO36), .W6(W6TO36), .W7(W7TO36), .W8(W8TO36), .W9(W9TO36), .W10(W10TO36), .W11(W11TO36), .W12(W12TO36), .W13(W13TO36), .W14(W14TO36), .W15(W15TO36), .W16(W16TO36), .W17(W17TO36), .W18(W18TO36), .W19(W19TO36), .W20(W20TO36), .W21(W21TO36), .W22(W22TO36), .W23(W23TO36), .W24(W24TO36), .W25(W25TO36), .W26(W26TO36), .W27(W27TO36), .W28(W28TO36), .W29(W29TO36), .W30(W30TO36), .W31(W31TO36), .W32(W32TO36), .W33(W33TO36), .W34(W34TO36), .W35(W35TO36), .W36(W36TO36), .W37(W37TO36), .W38(W38TO36), .W39(W39TO36), .W40(W40TO36), .W41(W41TO36), .W42(W42TO36), .W43(W43TO36), .W44(W44TO36), .W45(W45TO36), .W46(W46TO36), .W47(W47TO36), .W48(W48TO36), .W49(W49TO36), .W50(W50TO36), .W51(W51TO36), .W52(W52TO36), .W53(W53TO36), .W54(W54TO36), .W55(W55TO36), .W56(W56TO36), .W57(W57TO36), .W58(W58TO36), .W59(W59TO36), .W60(W60TO36), .W61(W61TO36), .W62(W62TO36), .W63(W63TO36), .W64(W64TO36)) neuron36(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out36));
neuron65in #(.BIAS(BIAS37), .W0(W0TO37), .W1(W1TO37), .W2(W2TO37), .W3(W3TO37), .W4(W4TO37), .W5(W5TO37), .W6(W6TO37), .W7(W7TO37), .W8(W8TO37), .W9(W9TO37), .W10(W10TO37), .W11(W11TO37), .W12(W12TO37), .W13(W13TO37), .W14(W14TO37), .W15(W15TO37), .W16(W16TO37), .W17(W17TO37), .W18(W18TO37), .W19(W19TO37), .W20(W20TO37), .W21(W21TO37), .W22(W22TO37), .W23(W23TO37), .W24(W24TO37), .W25(W25TO37), .W26(W26TO37), .W27(W27TO37), .W28(W28TO37), .W29(W29TO37), .W30(W30TO37), .W31(W31TO37), .W32(W32TO37), .W33(W33TO37), .W34(W34TO37), .W35(W35TO37), .W36(W36TO37), .W37(W37TO37), .W38(W38TO37), .W39(W39TO37), .W40(W40TO37), .W41(W41TO37), .W42(W42TO37), .W43(W43TO37), .W44(W44TO37), .W45(W45TO37), .W46(W46TO37), .W47(W47TO37), .W48(W48TO37), .W49(W49TO37), .W50(W50TO37), .W51(W51TO37), .W52(W52TO37), .W53(W53TO37), .W54(W54TO37), .W55(W55TO37), .W56(W56TO37), .W57(W57TO37), .W58(W58TO37), .W59(W59TO37), .W60(W60TO37), .W61(W61TO37), .W62(W62TO37), .W63(W63TO37), .W64(W64TO37)) neuron37(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out37));
neuron65in #(.BIAS(BIAS38), .W0(W0TO38), .W1(W1TO38), .W2(W2TO38), .W3(W3TO38), .W4(W4TO38), .W5(W5TO38), .W6(W6TO38), .W7(W7TO38), .W8(W8TO38), .W9(W9TO38), .W10(W10TO38), .W11(W11TO38), .W12(W12TO38), .W13(W13TO38), .W14(W14TO38), .W15(W15TO38), .W16(W16TO38), .W17(W17TO38), .W18(W18TO38), .W19(W19TO38), .W20(W20TO38), .W21(W21TO38), .W22(W22TO38), .W23(W23TO38), .W24(W24TO38), .W25(W25TO38), .W26(W26TO38), .W27(W27TO38), .W28(W28TO38), .W29(W29TO38), .W30(W30TO38), .W31(W31TO38), .W32(W32TO38), .W33(W33TO38), .W34(W34TO38), .W35(W35TO38), .W36(W36TO38), .W37(W37TO38), .W38(W38TO38), .W39(W39TO38), .W40(W40TO38), .W41(W41TO38), .W42(W42TO38), .W43(W43TO38), .W44(W44TO38), .W45(W45TO38), .W46(W46TO38), .W47(W47TO38), .W48(W48TO38), .W49(W49TO38), .W50(W50TO38), .W51(W51TO38), .W52(W52TO38), .W53(W53TO38), .W54(W54TO38), .W55(W55TO38), .W56(W56TO38), .W57(W57TO38), .W58(W58TO38), .W59(W59TO38), .W60(W60TO38), .W61(W61TO38), .W62(W62TO38), .W63(W63TO38), .W64(W64TO38)) neuron38(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out38));
neuron65in #(.BIAS(BIAS39), .W0(W0TO39), .W1(W1TO39), .W2(W2TO39), .W3(W3TO39), .W4(W4TO39), .W5(W5TO39), .W6(W6TO39), .W7(W7TO39), .W8(W8TO39), .W9(W9TO39), .W10(W10TO39), .W11(W11TO39), .W12(W12TO39), .W13(W13TO39), .W14(W14TO39), .W15(W15TO39), .W16(W16TO39), .W17(W17TO39), .W18(W18TO39), .W19(W19TO39), .W20(W20TO39), .W21(W21TO39), .W22(W22TO39), .W23(W23TO39), .W24(W24TO39), .W25(W25TO39), .W26(W26TO39), .W27(W27TO39), .W28(W28TO39), .W29(W29TO39), .W30(W30TO39), .W31(W31TO39), .W32(W32TO39), .W33(W33TO39), .W34(W34TO39), .W35(W35TO39), .W36(W36TO39), .W37(W37TO39), .W38(W38TO39), .W39(W39TO39), .W40(W40TO39), .W41(W41TO39), .W42(W42TO39), .W43(W43TO39), .W44(W44TO39), .W45(W45TO39), .W46(W46TO39), .W47(W47TO39), .W48(W48TO39), .W49(W49TO39), .W50(W50TO39), .W51(W51TO39), .W52(W52TO39), .W53(W53TO39), .W54(W54TO39), .W55(W55TO39), .W56(W56TO39), .W57(W57TO39), .W58(W58TO39), .W59(W59TO39), .W60(W60TO39), .W61(W61TO39), .W62(W62TO39), .W63(W63TO39), .W64(W64TO39)) neuron39(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out39));
neuron65in #(.BIAS(BIAS40), .W0(W0TO40), .W1(W1TO40), .W2(W2TO40), .W3(W3TO40), .W4(W4TO40), .W5(W5TO40), .W6(W6TO40), .W7(W7TO40), .W8(W8TO40), .W9(W9TO40), .W10(W10TO40), .W11(W11TO40), .W12(W12TO40), .W13(W13TO40), .W14(W14TO40), .W15(W15TO40), .W16(W16TO40), .W17(W17TO40), .W18(W18TO40), .W19(W19TO40), .W20(W20TO40), .W21(W21TO40), .W22(W22TO40), .W23(W23TO40), .W24(W24TO40), .W25(W25TO40), .W26(W26TO40), .W27(W27TO40), .W28(W28TO40), .W29(W29TO40), .W30(W30TO40), .W31(W31TO40), .W32(W32TO40), .W33(W33TO40), .W34(W34TO40), .W35(W35TO40), .W36(W36TO40), .W37(W37TO40), .W38(W38TO40), .W39(W39TO40), .W40(W40TO40), .W41(W41TO40), .W42(W42TO40), .W43(W43TO40), .W44(W44TO40), .W45(W45TO40), .W46(W46TO40), .W47(W47TO40), .W48(W48TO40), .W49(W49TO40), .W50(W50TO40), .W51(W51TO40), .W52(W52TO40), .W53(W53TO40), .W54(W54TO40), .W55(W55TO40), .W56(W56TO40), .W57(W57TO40), .W58(W58TO40), .W59(W59TO40), .W60(W60TO40), .W61(W61TO40), .W62(W62TO40), .W63(W63TO40), .W64(W64TO40)) neuron40(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out40));
neuron65in #(.BIAS(BIAS41), .W0(W0TO41), .W1(W1TO41), .W2(W2TO41), .W3(W3TO41), .W4(W4TO41), .W5(W5TO41), .W6(W6TO41), .W7(W7TO41), .W8(W8TO41), .W9(W9TO41), .W10(W10TO41), .W11(W11TO41), .W12(W12TO41), .W13(W13TO41), .W14(W14TO41), .W15(W15TO41), .W16(W16TO41), .W17(W17TO41), .W18(W18TO41), .W19(W19TO41), .W20(W20TO41), .W21(W21TO41), .W22(W22TO41), .W23(W23TO41), .W24(W24TO41), .W25(W25TO41), .W26(W26TO41), .W27(W27TO41), .W28(W28TO41), .W29(W29TO41), .W30(W30TO41), .W31(W31TO41), .W32(W32TO41), .W33(W33TO41), .W34(W34TO41), .W35(W35TO41), .W36(W36TO41), .W37(W37TO41), .W38(W38TO41), .W39(W39TO41), .W40(W40TO41), .W41(W41TO41), .W42(W42TO41), .W43(W43TO41), .W44(W44TO41), .W45(W45TO41), .W46(W46TO41), .W47(W47TO41), .W48(W48TO41), .W49(W49TO41), .W50(W50TO41), .W51(W51TO41), .W52(W52TO41), .W53(W53TO41), .W54(W54TO41), .W55(W55TO41), .W56(W56TO41), .W57(W57TO41), .W58(W58TO41), .W59(W59TO41), .W60(W60TO41), .W61(W61TO41), .W62(W62TO41), .W63(W63TO41), .W64(W64TO41)) neuron41(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out41));
neuron65in #(.BIAS(BIAS42), .W0(W0TO42), .W1(W1TO42), .W2(W2TO42), .W3(W3TO42), .W4(W4TO42), .W5(W5TO42), .W6(W6TO42), .W7(W7TO42), .W8(W8TO42), .W9(W9TO42), .W10(W10TO42), .W11(W11TO42), .W12(W12TO42), .W13(W13TO42), .W14(W14TO42), .W15(W15TO42), .W16(W16TO42), .W17(W17TO42), .W18(W18TO42), .W19(W19TO42), .W20(W20TO42), .W21(W21TO42), .W22(W22TO42), .W23(W23TO42), .W24(W24TO42), .W25(W25TO42), .W26(W26TO42), .W27(W27TO42), .W28(W28TO42), .W29(W29TO42), .W30(W30TO42), .W31(W31TO42), .W32(W32TO42), .W33(W33TO42), .W34(W34TO42), .W35(W35TO42), .W36(W36TO42), .W37(W37TO42), .W38(W38TO42), .W39(W39TO42), .W40(W40TO42), .W41(W41TO42), .W42(W42TO42), .W43(W43TO42), .W44(W44TO42), .W45(W45TO42), .W46(W46TO42), .W47(W47TO42), .W48(W48TO42), .W49(W49TO42), .W50(W50TO42), .W51(W51TO42), .W52(W52TO42), .W53(W53TO42), .W54(W54TO42), .W55(W55TO42), .W56(W56TO42), .W57(W57TO42), .W58(W58TO42), .W59(W59TO42), .W60(W60TO42), .W61(W61TO42), .W62(W62TO42), .W63(W63TO42), .W64(W64TO42)) neuron42(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out42));
neuron65in #(.BIAS(BIAS43), .W0(W0TO43), .W1(W1TO43), .W2(W2TO43), .W3(W3TO43), .W4(W4TO43), .W5(W5TO43), .W6(W6TO43), .W7(W7TO43), .W8(W8TO43), .W9(W9TO43), .W10(W10TO43), .W11(W11TO43), .W12(W12TO43), .W13(W13TO43), .W14(W14TO43), .W15(W15TO43), .W16(W16TO43), .W17(W17TO43), .W18(W18TO43), .W19(W19TO43), .W20(W20TO43), .W21(W21TO43), .W22(W22TO43), .W23(W23TO43), .W24(W24TO43), .W25(W25TO43), .W26(W26TO43), .W27(W27TO43), .W28(W28TO43), .W29(W29TO43), .W30(W30TO43), .W31(W31TO43), .W32(W32TO43), .W33(W33TO43), .W34(W34TO43), .W35(W35TO43), .W36(W36TO43), .W37(W37TO43), .W38(W38TO43), .W39(W39TO43), .W40(W40TO43), .W41(W41TO43), .W42(W42TO43), .W43(W43TO43), .W44(W44TO43), .W45(W45TO43), .W46(W46TO43), .W47(W47TO43), .W48(W48TO43), .W49(W49TO43), .W50(W50TO43), .W51(W51TO43), .W52(W52TO43), .W53(W53TO43), .W54(W54TO43), .W55(W55TO43), .W56(W56TO43), .W57(W57TO43), .W58(W58TO43), .W59(W59TO43), .W60(W60TO43), .W61(W61TO43), .W62(W62TO43), .W63(W63TO43), .W64(W64TO43)) neuron43(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out43));
neuron65in #(.BIAS(BIAS44), .W0(W0TO44), .W1(W1TO44), .W2(W2TO44), .W3(W3TO44), .W4(W4TO44), .W5(W5TO44), .W6(W6TO44), .W7(W7TO44), .W8(W8TO44), .W9(W9TO44), .W10(W10TO44), .W11(W11TO44), .W12(W12TO44), .W13(W13TO44), .W14(W14TO44), .W15(W15TO44), .W16(W16TO44), .W17(W17TO44), .W18(W18TO44), .W19(W19TO44), .W20(W20TO44), .W21(W21TO44), .W22(W22TO44), .W23(W23TO44), .W24(W24TO44), .W25(W25TO44), .W26(W26TO44), .W27(W27TO44), .W28(W28TO44), .W29(W29TO44), .W30(W30TO44), .W31(W31TO44), .W32(W32TO44), .W33(W33TO44), .W34(W34TO44), .W35(W35TO44), .W36(W36TO44), .W37(W37TO44), .W38(W38TO44), .W39(W39TO44), .W40(W40TO44), .W41(W41TO44), .W42(W42TO44), .W43(W43TO44), .W44(W44TO44), .W45(W45TO44), .W46(W46TO44), .W47(W47TO44), .W48(W48TO44), .W49(W49TO44), .W50(W50TO44), .W51(W51TO44), .W52(W52TO44), .W53(W53TO44), .W54(W54TO44), .W55(W55TO44), .W56(W56TO44), .W57(W57TO44), .W58(W58TO44), .W59(W59TO44), .W60(W60TO44), .W61(W61TO44), .W62(W62TO44), .W63(W63TO44), .W64(W64TO44)) neuron44(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out44));
neuron65in #(.BIAS(BIAS45), .W0(W0TO45), .W1(W1TO45), .W2(W2TO45), .W3(W3TO45), .W4(W4TO45), .W5(W5TO45), .W6(W6TO45), .W7(W7TO45), .W8(W8TO45), .W9(W9TO45), .W10(W10TO45), .W11(W11TO45), .W12(W12TO45), .W13(W13TO45), .W14(W14TO45), .W15(W15TO45), .W16(W16TO45), .W17(W17TO45), .W18(W18TO45), .W19(W19TO45), .W20(W20TO45), .W21(W21TO45), .W22(W22TO45), .W23(W23TO45), .W24(W24TO45), .W25(W25TO45), .W26(W26TO45), .W27(W27TO45), .W28(W28TO45), .W29(W29TO45), .W30(W30TO45), .W31(W31TO45), .W32(W32TO45), .W33(W33TO45), .W34(W34TO45), .W35(W35TO45), .W36(W36TO45), .W37(W37TO45), .W38(W38TO45), .W39(W39TO45), .W40(W40TO45), .W41(W41TO45), .W42(W42TO45), .W43(W43TO45), .W44(W44TO45), .W45(W45TO45), .W46(W46TO45), .W47(W47TO45), .W48(W48TO45), .W49(W49TO45), .W50(W50TO45), .W51(W51TO45), .W52(W52TO45), .W53(W53TO45), .W54(W54TO45), .W55(W55TO45), .W56(W56TO45), .W57(W57TO45), .W58(W58TO45), .W59(W59TO45), .W60(W60TO45), .W61(W61TO45), .W62(W62TO45), .W63(W63TO45), .W64(W64TO45)) neuron45(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out45));
neuron65in #(.BIAS(BIAS46), .W0(W0TO46), .W1(W1TO46), .W2(W2TO46), .W3(W3TO46), .W4(W4TO46), .W5(W5TO46), .W6(W6TO46), .W7(W7TO46), .W8(W8TO46), .W9(W9TO46), .W10(W10TO46), .W11(W11TO46), .W12(W12TO46), .W13(W13TO46), .W14(W14TO46), .W15(W15TO46), .W16(W16TO46), .W17(W17TO46), .W18(W18TO46), .W19(W19TO46), .W20(W20TO46), .W21(W21TO46), .W22(W22TO46), .W23(W23TO46), .W24(W24TO46), .W25(W25TO46), .W26(W26TO46), .W27(W27TO46), .W28(W28TO46), .W29(W29TO46), .W30(W30TO46), .W31(W31TO46), .W32(W32TO46), .W33(W33TO46), .W34(W34TO46), .W35(W35TO46), .W36(W36TO46), .W37(W37TO46), .W38(W38TO46), .W39(W39TO46), .W40(W40TO46), .W41(W41TO46), .W42(W42TO46), .W43(W43TO46), .W44(W44TO46), .W45(W45TO46), .W46(W46TO46), .W47(W47TO46), .W48(W48TO46), .W49(W49TO46), .W50(W50TO46), .W51(W51TO46), .W52(W52TO46), .W53(W53TO46), .W54(W54TO46), .W55(W55TO46), .W56(W56TO46), .W57(W57TO46), .W58(W58TO46), .W59(W59TO46), .W60(W60TO46), .W61(W61TO46), .W62(W62TO46), .W63(W63TO46), .W64(W64TO46)) neuron46(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out46));
neuron65in #(.BIAS(BIAS47), .W0(W0TO47), .W1(W1TO47), .W2(W2TO47), .W3(W3TO47), .W4(W4TO47), .W5(W5TO47), .W6(W6TO47), .W7(W7TO47), .W8(W8TO47), .W9(W9TO47), .W10(W10TO47), .W11(W11TO47), .W12(W12TO47), .W13(W13TO47), .W14(W14TO47), .W15(W15TO47), .W16(W16TO47), .W17(W17TO47), .W18(W18TO47), .W19(W19TO47), .W20(W20TO47), .W21(W21TO47), .W22(W22TO47), .W23(W23TO47), .W24(W24TO47), .W25(W25TO47), .W26(W26TO47), .W27(W27TO47), .W28(W28TO47), .W29(W29TO47), .W30(W30TO47), .W31(W31TO47), .W32(W32TO47), .W33(W33TO47), .W34(W34TO47), .W35(W35TO47), .W36(W36TO47), .W37(W37TO47), .W38(W38TO47), .W39(W39TO47), .W40(W40TO47), .W41(W41TO47), .W42(W42TO47), .W43(W43TO47), .W44(W44TO47), .W45(W45TO47), .W46(W46TO47), .W47(W47TO47), .W48(W48TO47), .W49(W49TO47), .W50(W50TO47), .W51(W51TO47), .W52(W52TO47), .W53(W53TO47), .W54(W54TO47), .W55(W55TO47), .W56(W56TO47), .W57(W57TO47), .W58(W58TO47), .W59(W59TO47), .W60(W60TO47), .W61(W61TO47), .W62(W62TO47), .W63(W63TO47), .W64(W64TO47)) neuron47(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out47));
neuron65in #(.BIAS(BIAS48), .W0(W0TO48), .W1(W1TO48), .W2(W2TO48), .W3(W3TO48), .W4(W4TO48), .W5(W5TO48), .W6(W6TO48), .W7(W7TO48), .W8(W8TO48), .W9(W9TO48), .W10(W10TO48), .W11(W11TO48), .W12(W12TO48), .W13(W13TO48), .W14(W14TO48), .W15(W15TO48), .W16(W16TO48), .W17(W17TO48), .W18(W18TO48), .W19(W19TO48), .W20(W20TO48), .W21(W21TO48), .W22(W22TO48), .W23(W23TO48), .W24(W24TO48), .W25(W25TO48), .W26(W26TO48), .W27(W27TO48), .W28(W28TO48), .W29(W29TO48), .W30(W30TO48), .W31(W31TO48), .W32(W32TO48), .W33(W33TO48), .W34(W34TO48), .W35(W35TO48), .W36(W36TO48), .W37(W37TO48), .W38(W38TO48), .W39(W39TO48), .W40(W40TO48), .W41(W41TO48), .W42(W42TO48), .W43(W43TO48), .W44(W44TO48), .W45(W45TO48), .W46(W46TO48), .W47(W47TO48), .W48(W48TO48), .W49(W49TO48), .W50(W50TO48), .W51(W51TO48), .W52(W52TO48), .W53(W53TO48), .W54(W54TO48), .W55(W55TO48), .W56(W56TO48), .W57(W57TO48), .W58(W58TO48), .W59(W59TO48), .W60(W60TO48), .W61(W61TO48), .W62(W62TO48), .W63(W63TO48), .W64(W64TO48)) neuron48(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out48));
neuron65in #(.BIAS(BIAS49), .W0(W0TO49), .W1(W1TO49), .W2(W2TO49), .W3(W3TO49), .W4(W4TO49), .W5(W5TO49), .W6(W6TO49), .W7(W7TO49), .W8(W8TO49), .W9(W9TO49), .W10(W10TO49), .W11(W11TO49), .W12(W12TO49), .W13(W13TO49), .W14(W14TO49), .W15(W15TO49), .W16(W16TO49), .W17(W17TO49), .W18(W18TO49), .W19(W19TO49), .W20(W20TO49), .W21(W21TO49), .W22(W22TO49), .W23(W23TO49), .W24(W24TO49), .W25(W25TO49), .W26(W26TO49), .W27(W27TO49), .W28(W28TO49), .W29(W29TO49), .W30(W30TO49), .W31(W31TO49), .W32(W32TO49), .W33(W33TO49), .W34(W34TO49), .W35(W35TO49), .W36(W36TO49), .W37(W37TO49), .W38(W38TO49), .W39(W39TO49), .W40(W40TO49), .W41(W41TO49), .W42(W42TO49), .W43(W43TO49), .W44(W44TO49), .W45(W45TO49), .W46(W46TO49), .W47(W47TO49), .W48(W48TO49), .W49(W49TO49), .W50(W50TO49), .W51(W51TO49), .W52(W52TO49), .W53(W53TO49), .W54(W54TO49), .W55(W55TO49), .W56(W56TO49), .W57(W57TO49), .W58(W58TO49), .W59(W59TO49), .W60(W60TO49), .W61(W61TO49), .W62(W62TO49), .W63(W63TO49), .W64(W64TO49)) neuron49(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out49));
neuron65in #(.BIAS(BIAS50), .W0(W0TO50), .W1(W1TO50), .W2(W2TO50), .W3(W3TO50), .W4(W4TO50), .W5(W5TO50), .W6(W6TO50), .W7(W7TO50), .W8(W8TO50), .W9(W9TO50), .W10(W10TO50), .W11(W11TO50), .W12(W12TO50), .W13(W13TO50), .W14(W14TO50), .W15(W15TO50), .W16(W16TO50), .W17(W17TO50), .W18(W18TO50), .W19(W19TO50), .W20(W20TO50), .W21(W21TO50), .W22(W22TO50), .W23(W23TO50), .W24(W24TO50), .W25(W25TO50), .W26(W26TO50), .W27(W27TO50), .W28(W28TO50), .W29(W29TO50), .W30(W30TO50), .W31(W31TO50), .W32(W32TO50), .W33(W33TO50), .W34(W34TO50), .W35(W35TO50), .W36(W36TO50), .W37(W37TO50), .W38(W38TO50), .W39(W39TO50), .W40(W40TO50), .W41(W41TO50), .W42(W42TO50), .W43(W43TO50), .W44(W44TO50), .W45(W45TO50), .W46(W46TO50), .W47(W47TO50), .W48(W48TO50), .W49(W49TO50), .W50(W50TO50), .W51(W51TO50), .W52(W52TO50), .W53(W53TO50), .W54(W54TO50), .W55(W55TO50), .W56(W56TO50), .W57(W57TO50), .W58(W58TO50), .W59(W59TO50), .W60(W60TO50), .W61(W61TO50), .W62(W62TO50), .W63(W63TO50), .W64(W64TO50)) neuron50(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out50));
neuron65in #(.BIAS(BIAS51), .W0(W0TO51), .W1(W1TO51), .W2(W2TO51), .W3(W3TO51), .W4(W4TO51), .W5(W5TO51), .W6(W6TO51), .W7(W7TO51), .W8(W8TO51), .W9(W9TO51), .W10(W10TO51), .W11(W11TO51), .W12(W12TO51), .W13(W13TO51), .W14(W14TO51), .W15(W15TO51), .W16(W16TO51), .W17(W17TO51), .W18(W18TO51), .W19(W19TO51), .W20(W20TO51), .W21(W21TO51), .W22(W22TO51), .W23(W23TO51), .W24(W24TO51), .W25(W25TO51), .W26(W26TO51), .W27(W27TO51), .W28(W28TO51), .W29(W29TO51), .W30(W30TO51), .W31(W31TO51), .W32(W32TO51), .W33(W33TO51), .W34(W34TO51), .W35(W35TO51), .W36(W36TO51), .W37(W37TO51), .W38(W38TO51), .W39(W39TO51), .W40(W40TO51), .W41(W41TO51), .W42(W42TO51), .W43(W43TO51), .W44(W44TO51), .W45(W45TO51), .W46(W46TO51), .W47(W47TO51), .W48(W48TO51), .W49(W49TO51), .W50(W50TO51), .W51(W51TO51), .W52(W52TO51), .W53(W53TO51), .W54(W54TO51), .W55(W55TO51), .W56(W56TO51), .W57(W57TO51), .W58(W58TO51), .W59(W59TO51), .W60(W60TO51), .W61(W61TO51), .W62(W62TO51), .W63(W63TO51), .W64(W64TO51)) neuron51(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out51));
neuron65in #(.BIAS(BIAS52), .W0(W0TO52), .W1(W1TO52), .W2(W2TO52), .W3(W3TO52), .W4(W4TO52), .W5(W5TO52), .W6(W6TO52), .W7(W7TO52), .W8(W8TO52), .W9(W9TO52), .W10(W10TO52), .W11(W11TO52), .W12(W12TO52), .W13(W13TO52), .W14(W14TO52), .W15(W15TO52), .W16(W16TO52), .W17(W17TO52), .W18(W18TO52), .W19(W19TO52), .W20(W20TO52), .W21(W21TO52), .W22(W22TO52), .W23(W23TO52), .W24(W24TO52), .W25(W25TO52), .W26(W26TO52), .W27(W27TO52), .W28(W28TO52), .W29(W29TO52), .W30(W30TO52), .W31(W31TO52), .W32(W32TO52), .W33(W33TO52), .W34(W34TO52), .W35(W35TO52), .W36(W36TO52), .W37(W37TO52), .W38(W38TO52), .W39(W39TO52), .W40(W40TO52), .W41(W41TO52), .W42(W42TO52), .W43(W43TO52), .W44(W44TO52), .W45(W45TO52), .W46(W46TO52), .W47(W47TO52), .W48(W48TO52), .W49(W49TO52), .W50(W50TO52), .W51(W51TO52), .W52(W52TO52), .W53(W53TO52), .W54(W54TO52), .W55(W55TO52), .W56(W56TO52), .W57(W57TO52), .W58(W58TO52), .W59(W59TO52), .W60(W60TO52), .W61(W61TO52), .W62(W62TO52), .W63(W63TO52), .W64(W64TO52)) neuron52(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out52));
neuron65in #(.BIAS(BIAS53), .W0(W0TO53), .W1(W1TO53), .W2(W2TO53), .W3(W3TO53), .W4(W4TO53), .W5(W5TO53), .W6(W6TO53), .W7(W7TO53), .W8(W8TO53), .W9(W9TO53), .W10(W10TO53), .W11(W11TO53), .W12(W12TO53), .W13(W13TO53), .W14(W14TO53), .W15(W15TO53), .W16(W16TO53), .W17(W17TO53), .W18(W18TO53), .W19(W19TO53), .W20(W20TO53), .W21(W21TO53), .W22(W22TO53), .W23(W23TO53), .W24(W24TO53), .W25(W25TO53), .W26(W26TO53), .W27(W27TO53), .W28(W28TO53), .W29(W29TO53), .W30(W30TO53), .W31(W31TO53), .W32(W32TO53), .W33(W33TO53), .W34(W34TO53), .W35(W35TO53), .W36(W36TO53), .W37(W37TO53), .W38(W38TO53), .W39(W39TO53), .W40(W40TO53), .W41(W41TO53), .W42(W42TO53), .W43(W43TO53), .W44(W44TO53), .W45(W45TO53), .W46(W46TO53), .W47(W47TO53), .W48(W48TO53), .W49(W49TO53), .W50(W50TO53), .W51(W51TO53), .W52(W52TO53), .W53(W53TO53), .W54(W54TO53), .W55(W55TO53), .W56(W56TO53), .W57(W57TO53), .W58(W58TO53), .W59(W59TO53), .W60(W60TO53), .W61(W61TO53), .W62(W62TO53), .W63(W63TO53), .W64(W64TO53)) neuron53(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out53));
neuron65in #(.BIAS(BIAS54), .W0(W0TO54), .W1(W1TO54), .W2(W2TO54), .W3(W3TO54), .W4(W4TO54), .W5(W5TO54), .W6(W6TO54), .W7(W7TO54), .W8(W8TO54), .W9(W9TO54), .W10(W10TO54), .W11(W11TO54), .W12(W12TO54), .W13(W13TO54), .W14(W14TO54), .W15(W15TO54), .W16(W16TO54), .W17(W17TO54), .W18(W18TO54), .W19(W19TO54), .W20(W20TO54), .W21(W21TO54), .W22(W22TO54), .W23(W23TO54), .W24(W24TO54), .W25(W25TO54), .W26(W26TO54), .W27(W27TO54), .W28(W28TO54), .W29(W29TO54), .W30(W30TO54), .W31(W31TO54), .W32(W32TO54), .W33(W33TO54), .W34(W34TO54), .W35(W35TO54), .W36(W36TO54), .W37(W37TO54), .W38(W38TO54), .W39(W39TO54), .W40(W40TO54), .W41(W41TO54), .W42(W42TO54), .W43(W43TO54), .W44(W44TO54), .W45(W45TO54), .W46(W46TO54), .W47(W47TO54), .W48(W48TO54), .W49(W49TO54), .W50(W50TO54), .W51(W51TO54), .W52(W52TO54), .W53(W53TO54), .W54(W54TO54), .W55(W55TO54), .W56(W56TO54), .W57(W57TO54), .W58(W58TO54), .W59(W59TO54), .W60(W60TO54), .W61(W61TO54), .W62(W62TO54), .W63(W63TO54), .W64(W64TO54)) neuron54(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out54));
neuron65in #(.BIAS(BIAS55), .W0(W0TO55), .W1(W1TO55), .W2(W2TO55), .W3(W3TO55), .W4(W4TO55), .W5(W5TO55), .W6(W6TO55), .W7(W7TO55), .W8(W8TO55), .W9(W9TO55), .W10(W10TO55), .W11(W11TO55), .W12(W12TO55), .W13(W13TO55), .W14(W14TO55), .W15(W15TO55), .W16(W16TO55), .W17(W17TO55), .W18(W18TO55), .W19(W19TO55), .W20(W20TO55), .W21(W21TO55), .W22(W22TO55), .W23(W23TO55), .W24(W24TO55), .W25(W25TO55), .W26(W26TO55), .W27(W27TO55), .W28(W28TO55), .W29(W29TO55), .W30(W30TO55), .W31(W31TO55), .W32(W32TO55), .W33(W33TO55), .W34(W34TO55), .W35(W35TO55), .W36(W36TO55), .W37(W37TO55), .W38(W38TO55), .W39(W39TO55), .W40(W40TO55), .W41(W41TO55), .W42(W42TO55), .W43(W43TO55), .W44(W44TO55), .W45(W45TO55), .W46(W46TO55), .W47(W47TO55), .W48(W48TO55), .W49(W49TO55), .W50(W50TO55), .W51(W51TO55), .W52(W52TO55), .W53(W53TO55), .W54(W54TO55), .W55(W55TO55), .W56(W56TO55), .W57(W57TO55), .W58(W58TO55), .W59(W59TO55), .W60(W60TO55), .W61(W61TO55), .W62(W62TO55), .W63(W63TO55), .W64(W64TO55)) neuron55(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out55));
neuron65in #(.BIAS(BIAS56), .W0(W0TO56), .W1(W1TO56), .W2(W2TO56), .W3(W3TO56), .W4(W4TO56), .W5(W5TO56), .W6(W6TO56), .W7(W7TO56), .W8(W8TO56), .W9(W9TO56), .W10(W10TO56), .W11(W11TO56), .W12(W12TO56), .W13(W13TO56), .W14(W14TO56), .W15(W15TO56), .W16(W16TO56), .W17(W17TO56), .W18(W18TO56), .W19(W19TO56), .W20(W20TO56), .W21(W21TO56), .W22(W22TO56), .W23(W23TO56), .W24(W24TO56), .W25(W25TO56), .W26(W26TO56), .W27(W27TO56), .W28(W28TO56), .W29(W29TO56), .W30(W30TO56), .W31(W31TO56), .W32(W32TO56), .W33(W33TO56), .W34(W34TO56), .W35(W35TO56), .W36(W36TO56), .W37(W37TO56), .W38(W38TO56), .W39(W39TO56), .W40(W40TO56), .W41(W41TO56), .W42(W42TO56), .W43(W43TO56), .W44(W44TO56), .W45(W45TO56), .W46(W46TO56), .W47(W47TO56), .W48(W48TO56), .W49(W49TO56), .W50(W50TO56), .W51(W51TO56), .W52(W52TO56), .W53(W53TO56), .W54(W54TO56), .W55(W55TO56), .W56(W56TO56), .W57(W57TO56), .W58(W58TO56), .W59(W59TO56), .W60(W60TO56), .W61(W61TO56), .W62(W62TO56), .W63(W63TO56), .W64(W64TO56)) neuron56(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out56));
neuron65in #(.BIAS(BIAS57), .W0(W0TO57), .W1(W1TO57), .W2(W2TO57), .W3(W3TO57), .W4(W4TO57), .W5(W5TO57), .W6(W6TO57), .W7(W7TO57), .W8(W8TO57), .W9(W9TO57), .W10(W10TO57), .W11(W11TO57), .W12(W12TO57), .W13(W13TO57), .W14(W14TO57), .W15(W15TO57), .W16(W16TO57), .W17(W17TO57), .W18(W18TO57), .W19(W19TO57), .W20(W20TO57), .W21(W21TO57), .W22(W22TO57), .W23(W23TO57), .W24(W24TO57), .W25(W25TO57), .W26(W26TO57), .W27(W27TO57), .W28(W28TO57), .W29(W29TO57), .W30(W30TO57), .W31(W31TO57), .W32(W32TO57), .W33(W33TO57), .W34(W34TO57), .W35(W35TO57), .W36(W36TO57), .W37(W37TO57), .W38(W38TO57), .W39(W39TO57), .W40(W40TO57), .W41(W41TO57), .W42(W42TO57), .W43(W43TO57), .W44(W44TO57), .W45(W45TO57), .W46(W46TO57), .W47(W47TO57), .W48(W48TO57), .W49(W49TO57), .W50(W50TO57), .W51(W51TO57), .W52(W52TO57), .W53(W53TO57), .W54(W54TO57), .W55(W55TO57), .W56(W56TO57), .W57(W57TO57), .W58(W58TO57), .W59(W59TO57), .W60(W60TO57), .W61(W61TO57), .W62(W62TO57), .W63(W63TO57), .W64(W64TO57)) neuron57(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out57));
neuron65in #(.BIAS(BIAS58), .W0(W0TO58), .W1(W1TO58), .W2(W2TO58), .W3(W3TO58), .W4(W4TO58), .W5(W5TO58), .W6(W6TO58), .W7(W7TO58), .W8(W8TO58), .W9(W9TO58), .W10(W10TO58), .W11(W11TO58), .W12(W12TO58), .W13(W13TO58), .W14(W14TO58), .W15(W15TO58), .W16(W16TO58), .W17(W17TO58), .W18(W18TO58), .W19(W19TO58), .W20(W20TO58), .W21(W21TO58), .W22(W22TO58), .W23(W23TO58), .W24(W24TO58), .W25(W25TO58), .W26(W26TO58), .W27(W27TO58), .W28(W28TO58), .W29(W29TO58), .W30(W30TO58), .W31(W31TO58), .W32(W32TO58), .W33(W33TO58), .W34(W34TO58), .W35(W35TO58), .W36(W36TO58), .W37(W37TO58), .W38(W38TO58), .W39(W39TO58), .W40(W40TO58), .W41(W41TO58), .W42(W42TO58), .W43(W43TO58), .W44(W44TO58), .W45(W45TO58), .W46(W46TO58), .W47(W47TO58), .W48(W48TO58), .W49(W49TO58), .W50(W50TO58), .W51(W51TO58), .W52(W52TO58), .W53(W53TO58), .W54(W54TO58), .W55(W55TO58), .W56(W56TO58), .W57(W57TO58), .W58(W58TO58), .W59(W59TO58), .W60(W60TO58), .W61(W61TO58), .W62(W62TO58), .W63(W63TO58), .W64(W64TO58)) neuron58(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out58));
neuron65in #(.BIAS(BIAS59), .W0(W0TO59), .W1(W1TO59), .W2(W2TO59), .W3(W3TO59), .W4(W4TO59), .W5(W5TO59), .W6(W6TO59), .W7(W7TO59), .W8(W8TO59), .W9(W9TO59), .W10(W10TO59), .W11(W11TO59), .W12(W12TO59), .W13(W13TO59), .W14(W14TO59), .W15(W15TO59), .W16(W16TO59), .W17(W17TO59), .W18(W18TO59), .W19(W19TO59), .W20(W20TO59), .W21(W21TO59), .W22(W22TO59), .W23(W23TO59), .W24(W24TO59), .W25(W25TO59), .W26(W26TO59), .W27(W27TO59), .W28(W28TO59), .W29(W29TO59), .W30(W30TO59), .W31(W31TO59), .W32(W32TO59), .W33(W33TO59), .W34(W34TO59), .W35(W35TO59), .W36(W36TO59), .W37(W37TO59), .W38(W38TO59), .W39(W39TO59), .W40(W40TO59), .W41(W41TO59), .W42(W42TO59), .W43(W43TO59), .W44(W44TO59), .W45(W45TO59), .W46(W46TO59), .W47(W47TO59), .W48(W48TO59), .W49(W49TO59), .W50(W50TO59), .W51(W51TO59), .W52(W52TO59), .W53(W53TO59), .W54(W54TO59), .W55(W55TO59), .W56(W56TO59), .W57(W57TO59), .W58(W58TO59), .W59(W59TO59), .W60(W60TO59), .W61(W61TO59), .W62(W62TO59), .W63(W63TO59), .W64(W64TO59)) neuron59(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out59));
neuron65in #(.BIAS(BIAS60), .W0(W0TO60), .W1(W1TO60), .W2(W2TO60), .W3(W3TO60), .W4(W4TO60), .W5(W5TO60), .W6(W6TO60), .W7(W7TO60), .W8(W8TO60), .W9(W9TO60), .W10(W10TO60), .W11(W11TO60), .W12(W12TO60), .W13(W13TO60), .W14(W14TO60), .W15(W15TO60), .W16(W16TO60), .W17(W17TO60), .W18(W18TO60), .W19(W19TO60), .W20(W20TO60), .W21(W21TO60), .W22(W22TO60), .W23(W23TO60), .W24(W24TO60), .W25(W25TO60), .W26(W26TO60), .W27(W27TO60), .W28(W28TO60), .W29(W29TO60), .W30(W30TO60), .W31(W31TO60), .W32(W32TO60), .W33(W33TO60), .W34(W34TO60), .W35(W35TO60), .W36(W36TO60), .W37(W37TO60), .W38(W38TO60), .W39(W39TO60), .W40(W40TO60), .W41(W41TO60), .W42(W42TO60), .W43(W43TO60), .W44(W44TO60), .W45(W45TO60), .W46(W46TO60), .W47(W47TO60), .W48(W48TO60), .W49(W49TO60), .W50(W50TO60), .W51(W51TO60), .W52(W52TO60), .W53(W53TO60), .W54(W54TO60), .W55(W55TO60), .W56(W56TO60), .W57(W57TO60), .W58(W58TO60), .W59(W59TO60), .W60(W60TO60), .W61(W61TO60), .W62(W62TO60), .W63(W63TO60), .W64(W64TO60)) neuron60(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out60));
neuron65in #(.BIAS(BIAS61), .W0(W0TO61), .W1(W1TO61), .W2(W2TO61), .W3(W3TO61), .W4(W4TO61), .W5(W5TO61), .W6(W6TO61), .W7(W7TO61), .W8(W8TO61), .W9(W9TO61), .W10(W10TO61), .W11(W11TO61), .W12(W12TO61), .W13(W13TO61), .W14(W14TO61), .W15(W15TO61), .W16(W16TO61), .W17(W17TO61), .W18(W18TO61), .W19(W19TO61), .W20(W20TO61), .W21(W21TO61), .W22(W22TO61), .W23(W23TO61), .W24(W24TO61), .W25(W25TO61), .W26(W26TO61), .W27(W27TO61), .W28(W28TO61), .W29(W29TO61), .W30(W30TO61), .W31(W31TO61), .W32(W32TO61), .W33(W33TO61), .W34(W34TO61), .W35(W35TO61), .W36(W36TO61), .W37(W37TO61), .W38(W38TO61), .W39(W39TO61), .W40(W40TO61), .W41(W41TO61), .W42(W42TO61), .W43(W43TO61), .W44(W44TO61), .W45(W45TO61), .W46(W46TO61), .W47(W47TO61), .W48(W48TO61), .W49(W49TO61), .W50(W50TO61), .W51(W51TO61), .W52(W52TO61), .W53(W53TO61), .W54(W54TO61), .W55(W55TO61), .W56(W56TO61), .W57(W57TO61), .W58(W58TO61), .W59(W59TO61), .W60(W60TO61), .W61(W61TO61), .W62(W62TO61), .W63(W63TO61), .W64(W64TO61)) neuron61(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out61));
neuron65in #(.BIAS(BIAS62), .W0(W0TO62), .W1(W1TO62), .W2(W2TO62), .W3(W3TO62), .W4(W4TO62), .W5(W5TO62), .W6(W6TO62), .W7(W7TO62), .W8(W8TO62), .W9(W9TO62), .W10(W10TO62), .W11(W11TO62), .W12(W12TO62), .W13(W13TO62), .W14(W14TO62), .W15(W15TO62), .W16(W16TO62), .W17(W17TO62), .W18(W18TO62), .W19(W19TO62), .W20(W20TO62), .W21(W21TO62), .W22(W22TO62), .W23(W23TO62), .W24(W24TO62), .W25(W25TO62), .W26(W26TO62), .W27(W27TO62), .W28(W28TO62), .W29(W29TO62), .W30(W30TO62), .W31(W31TO62), .W32(W32TO62), .W33(W33TO62), .W34(W34TO62), .W35(W35TO62), .W36(W36TO62), .W37(W37TO62), .W38(W38TO62), .W39(W39TO62), .W40(W40TO62), .W41(W41TO62), .W42(W42TO62), .W43(W43TO62), .W44(W44TO62), .W45(W45TO62), .W46(W46TO62), .W47(W47TO62), .W48(W48TO62), .W49(W49TO62), .W50(W50TO62), .W51(W51TO62), .W52(W52TO62), .W53(W53TO62), .W54(W54TO62), .W55(W55TO62), .W56(W56TO62), .W57(W57TO62), .W58(W58TO62), .W59(W59TO62), .W60(W60TO62), .W61(W61TO62), .W62(W62TO62), .W63(W63TO62), .W64(W64TO62)) neuron62(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out62));
neuron65in #(.BIAS(BIAS63), .W0(W0TO63), .W1(W1TO63), .W2(W2TO63), .W3(W3TO63), .W4(W4TO63), .W5(W5TO63), .W6(W6TO63), .W7(W7TO63), .W8(W8TO63), .W9(W9TO63), .W10(W10TO63), .W11(W11TO63), .W12(W12TO63), .W13(W13TO63), .W14(W14TO63), .W15(W15TO63), .W16(W16TO63), .W17(W17TO63), .W18(W18TO63), .W19(W19TO63), .W20(W20TO63), .W21(W21TO63), .W22(W22TO63), .W23(W23TO63), .W24(W24TO63), .W25(W25TO63), .W26(W26TO63), .W27(W27TO63), .W28(W28TO63), .W29(W29TO63), .W30(W30TO63), .W31(W31TO63), .W32(W32TO63), .W33(W33TO63), .W34(W34TO63), .W35(W35TO63), .W36(W36TO63), .W37(W37TO63), .W38(W38TO63), .W39(W39TO63), .W40(W40TO63), .W41(W41TO63), .W42(W42TO63), .W43(W43TO63), .W44(W44TO63), .W45(W45TO63), .W46(W46TO63), .W47(W47TO63), .W48(W48TO63), .W49(W49TO63), .W50(W50TO63), .W51(W51TO63), .W52(W52TO63), .W53(W53TO63), .W54(W54TO63), .W55(W55TO63), .W56(W56TO63), .W57(W57TO63), .W58(W58TO63), .W59(W59TO63), .W60(W60TO63), .W61(W61TO63), .W62(W62TO63), .W63(W63TO63), .W64(W64TO63)) neuron63(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out63));

endmodule

module layer64in1out(clk, rst, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, out0);

parameter signed BIAS0 = 0;
parameter signed W0TO0 = 0;
parameter signed W1TO0 = 0;
parameter signed W2TO0 = 0;
parameter signed W3TO0 = 0;
parameter signed W4TO0 = 0;
parameter signed W5TO0 = 0;
parameter signed W6TO0 = 0;
parameter signed W7TO0 = 0;
parameter signed W8TO0 = 0;
parameter signed W9TO0 = 0;
parameter signed W10TO0 = 0;
parameter signed W11TO0 = 0;
parameter signed W12TO0 = 0;
parameter signed W13TO0 = 0;
parameter signed W14TO0 = 0;
parameter signed W15TO0 = 0;
parameter signed W16TO0 = 0;
parameter signed W17TO0 = 0;
parameter signed W18TO0 = 0;
parameter signed W19TO0 = 0;
parameter signed W20TO0 = 0;
parameter signed W21TO0 = 0;
parameter signed W22TO0 = 0;
parameter signed W23TO0 = 0;
parameter signed W24TO0 = 0;
parameter signed W25TO0 = 0;
parameter signed W26TO0 = 0;
parameter signed W27TO0 = 0;
parameter signed W28TO0 = 0;
parameter signed W29TO0 = 0;
parameter signed W30TO0 = 0;
parameter signed W31TO0 = 0;
parameter signed W32TO0 = 0;
parameter signed W33TO0 = 0;
parameter signed W34TO0 = 0;
parameter signed W35TO0 = 0;
parameter signed W36TO0 = 0;
parameter signed W37TO0 = 0;
parameter signed W38TO0 = 0;
parameter signed W39TO0 = 0;
parameter signed W40TO0 = 0;
parameter signed W41TO0 = 0;
parameter signed W42TO0 = 0;
parameter signed W43TO0 = 0;
parameter signed W44TO0 = 0;
parameter signed W45TO0 = 0;
parameter signed W46TO0 = 0;
parameter signed W47TO0 = 0;
parameter signed W48TO0 = 0;
parameter signed W49TO0 = 0;
parameter signed W50TO0 = 0;
parameter signed W51TO0 = 0;
parameter signed W52TO0 = 0;
parameter signed W53TO0 = 0;
parameter signed W54TO0 = 0;
parameter signed W55TO0 = 0;
parameter signed W56TO0 = 0;
parameter signed W57TO0 = 0;
parameter signed W58TO0 = 0;
parameter signed W59TO0 = 0;
parameter signed W60TO0 = 0;
parameter signed W61TO0 = 0;
parameter signed W62TO0 = 0;
parameter signed W63TO0 = 0;

input wire clk;
input wire rst;

input signed [15:0] in0;
input signed [15:0] in1;
input signed [15:0] in2;
input signed [15:0] in3;
input signed [15:0] in4;
input signed [15:0] in5;
input signed [15:0] in6;
input signed [15:0] in7;
input signed [15:0] in8;
input signed [15:0] in9;
input signed [15:0] in10;
input signed [15:0] in11;
input signed [15:0] in12;
input signed [15:0] in13;
input signed [15:0] in14;
input signed [15:0] in15;
input signed [15:0] in16;
input signed [15:0] in17;
input signed [15:0] in18;
input signed [15:0] in19;
input signed [15:0] in20;
input signed [15:0] in21;
input signed [15:0] in22;
input signed [15:0] in23;
input signed [15:0] in24;
input signed [15:0] in25;
input signed [15:0] in26;
input signed [15:0] in27;
input signed [15:0] in28;
input signed [15:0] in29;
input signed [15:0] in30;
input signed [15:0] in31;
input signed [15:0] in32;
input signed [15:0] in33;
input signed [15:0] in34;
input signed [15:0] in35;
input signed [15:0] in36;
input signed [15:0] in37;
input signed [15:0] in38;
input signed [15:0] in39;
input signed [15:0] in40;
input signed [15:0] in41;
input signed [15:0] in42;
input signed [15:0] in43;
input signed [15:0] in44;
input signed [15:0] in45;
input signed [15:0] in46;
input signed [15:0] in47;
input signed [15:0] in48;
input signed [15:0] in49;
input signed [15:0] in50;
input signed [15:0] in51;
input signed [15:0] in52;
input signed [15:0] in53;
input signed [15:0] in54;
input signed [15:0] in55;
input signed [15:0] in56;
input signed [15:0] in57;
input signed [15:0] in58;
input signed [15:0] in59;
input signed [15:0] in60;
input signed [15:0] in61;
input signed [15:0] in62;
input signed [15:0] in63;

output signed [15:0] out0;

neuron64in #(.BIAS(BIAS0), .W0(W0TO0), .W1(W1TO0), .W2(W2TO0), .W3(W3TO0), .W4(W4TO0), .W5(W5TO0), .W6(W6TO0), .W7(W7TO0), .W8(W8TO0), .W9(W9TO0), .W10(W10TO0), .W11(W11TO0), .W12(W12TO0), .W13(W13TO0), .W14(W14TO0), .W15(W15TO0), .W16(W16TO0), .W17(W17TO0), .W18(W18TO0), .W19(W19TO0), .W20(W20TO0), .W21(W21TO0), .W22(W22TO0), .W23(W23TO0), .W24(W24TO0), .W25(W25TO0), .W26(W26TO0), .W27(W27TO0), .W28(W28TO0), .W29(W29TO0), .W30(W30TO0), .W31(W31TO0), .W32(W32TO0), .W33(W33TO0), .W34(W34TO0), .W35(W35TO0), .W36(W36TO0), .W37(W37TO0), .W38(W38TO0), .W39(W39TO0), .W40(W40TO0), .W41(W41TO0), .W42(W42TO0), .W43(W43TO0), .W44(W44TO0), .W45(W45TO0), .W46(W46TO0), .W47(W47TO0), .W48(W48TO0), .W49(W49TO0), .W50(W50TO0), .W51(W51TO0), .W52(W52TO0), .W53(W53TO0), .W54(W54TO0), .W55(W55TO0), .W56(W56TO0), .W57(W57TO0), .W58(W58TO0), .W59(W59TO0), .W60(W60TO0), .W61(W61TO0), .W62(W62TO0), .W63(W63TO0)) neuron0(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out0));

endmodule

module network(clk, rst, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, out0);

input wire clk;
input wire rst;

input signed [15:0] in0;
input signed [15:0] in1;
input signed [15:0] in2;
input signed [15:0] in3;
input signed [15:0] in4;
input signed [15:0] in5;
input signed [15:0] in6;
input signed [15:0] in7;
input signed [15:0] in8;
input signed [15:0] in9;
input signed [15:0] in10;
input signed [15:0] in11;
input signed [15:0] in12;
input signed [15:0] in13;
input signed [15:0] in14;
input signed [15:0] in15;
input signed [15:0] in16;
input signed [15:0] in17;
input signed [15:0] in18;
input signed [15:0] in19;
input signed [15:0] in20;
input signed [15:0] in21;
input signed [15:0] in22;
input signed [15:0] in23;
input signed [15:0] in24;
input signed [15:0] in25;
input signed [15:0] in26;
input signed [15:0] in27;
input signed [15:0] in28;
input signed [15:0] in29;
input signed [15:0] in30;
input signed [15:0] in31;
input signed [15:0] in32;
input signed [15:0] in33;
input signed [15:0] in34;
input signed [15:0] in35;
input signed [15:0] in36;
input signed [15:0] in37;
input signed [15:0] in38;
input signed [15:0] in39;
input signed [15:0] in40;
input signed [15:0] in41;
input signed [15:0] in42;
input signed [15:0] in43;
input signed [15:0] in44;
input signed [15:0] in45;
input signed [15:0] in46;
input signed [15:0] in47;
input signed [15:0] in48;
input signed [15:0] in49;
input signed [15:0] in50;
input signed [15:0] in51;
input signed [15:0] in52;
input signed [15:0] in53;
input signed [15:0] in54;
input signed [15:0] in55;
input signed [15:0] in56;
input signed [15:0] in57;
input signed [15:0] in58;
input signed [15:0] in59;
input signed [15:0] in60;
input signed [15:0] in61;
input signed [15:0] in62;
input signed [15:0] in63;
input signed [15:0] in64;

output signed [15:0] out0;

wire[15:0] con0[0:63];

layer65in64out #(.BIAS0(-475), .BIAS1(-682), .BIAS2(-443), .BIAS3(-80), .BIAS4(-357), .BIAS5(37), .BIAS6(-475), .BIAS7(952), .BIAS8(466), .BIAS9(-768), .BIAS10(-226), .BIAS11(257), .BIAS12(-749), .BIAS13(967), .BIAS14(-113), .BIAS15(579), .BIAS16(588), .BIAS17(-276), .BIAS18(-167), .BIAS19(169), .BIAS20(520), .BIAS21(-623), .BIAS22(-423), .BIAS23(340), .BIAS24(0), .BIAS25(-642), .BIAS26(-173), .BIAS27(-601), .BIAS28(63), .BIAS29(665), .BIAS30(-628), .BIAS31(915), .BIAS32(-148), .BIAS33(8), .BIAS34(21), .BIAS35(-967), .BIAS36(463), .BIAS37(987), .BIAS38(-673), .BIAS39(-746), .BIAS40(-249), .BIAS41(386), .BIAS42(-993), .BIAS43(-261), .BIAS44(-882), .BIAS45(579), .BIAS46(-299), .BIAS47(405), .BIAS48(-17), .BIAS49(946), .BIAS50(672), .BIAS51(220), .BIAS52(129), .BIAS53(995), .BIAS54(-490), .BIAS55(-970), .BIAS56(-821), .BIAS57(878), .BIAS58(947), .BIAS59(-16), .BIAS60(-317), .BIAS61(446), .BIAS62(-977), .BIAS63(520), .W0TO0(343), .W0TO1(-618), .W0TO2(333), .W0TO3(822), .W0TO4(-675), .W0TO5(821), .W0TO6(-350), .W0TO7(401), .W0TO8(-468), .W0TO9(38), .W0TO10(-644), .W0TO11(-63), .W0TO12(-101), .W0TO13(-207), .W0TO14(584), .W0TO15(-12), .W0TO16(448), .W0TO17(586), .W0TO18(-296), .W0TO19(819), .W0TO20(426), .W0TO21(794), .W0TO22(-159), .W0TO23(-64), .W0TO24(808), .W0TO25(267), .W0TO26(66), .W0TO27(-524), .W0TO28(893), .W0TO29(119), .W0TO30(515), .W0TO31(-527), .W0TO32(-139), .W0TO33(-211), .W0TO34(21), .W0TO35(-748), .W0TO36(367), .W0TO37(-944), .W0TO38(-531), .W0TO39(473), .W0TO40(868), .W0TO41(227), .W0TO42(-184), .W0TO43(708), .W0TO44(986), .W0TO45(-408), .W0TO46(-219), .W0TO47(398), .W0TO48(-285), .W0TO49(-935), .W0TO50(-301), .W0TO51(-29), .W0TO52(-903), .W0TO53(830), .W0TO54(451), .W0TO55(545), .W0TO56(-806), .W0TO57(-925), .W0TO58(-479), .W0TO59(-748), .W0TO60(-523), .W0TO61(364), .W0TO62(-37), .W0TO63(873), .W1TO0(163), .W1TO1(-627), .W1TO2(-625), .W1TO3(-322), .W1TO4(-133), .W1TO5(-845), .W1TO6(272), .W1TO7(-882), .W1TO8(447), .W1TO9(320), .W1TO10(-981), .W1TO11(526), .W1TO12(-322), .W1TO13(552), .W1TO14(-327), .W1TO15(161), .W1TO16(-655), .W1TO17(692), .W1TO18(-457), .W1TO19(489), .W1TO20(127), .W1TO21(800), .W1TO22(97), .W1TO23(-949), .W1TO24(-838), .W1TO25(911), .W1TO26(-87), .W1TO27(-704), .W1TO28(350), .W1TO29(247), .W1TO30(100), .W1TO31(812), .W1TO32(797), .W1TO33(-474), .W1TO34(438), .W1TO35(-29), .W1TO36(-437), .W1TO37(-882), .W1TO38(-589), .W1TO39(280), .W1TO40(-427), .W1TO41(-114), .W1TO42(-307), .W1TO43(0), .W1TO44(310), .W1TO45(899), .W1TO46(-933), .W1TO47(113), .W1TO48(282), .W1TO49(-682), .W1TO50(453), .W1TO51(-242), .W1TO52(23), .W1TO53(156), .W1TO54(691), .W1TO55(404), .W1TO56(258), .W1TO57(-896), .W1TO58(-907), .W1TO59(58), .W1TO60(566), .W1TO61(406), .W1TO62(-606), .W1TO63(-456), .W2TO0(-568), .W2TO1(-182), .W2TO2(311), .W2TO3(-458), .W2TO4(-438), .W2TO5(564), .W2TO6(704), .W2TO7(95), .W2TO8(448), .W2TO9(-133), .W2TO10(641), .W2TO11(649), .W2TO12(-966), .W2TO13(466), .W2TO14(434), .W2TO15(439), .W2TO16(572), .W2TO17(874), .W2TO18(316), .W2TO19(-624), .W2TO20(376), .W2TO21(981), .W2TO22(829), .W2TO23(730), .W2TO24(-906), .W2TO25(-983), .W2TO26(499), .W2TO27(467), .W2TO28(417), .W2TO29(-685), .W2TO30(-762), .W2TO31(-678), .W2TO32(646), .W2TO33(-192), .W2TO34(-641), .W2TO35(263), .W2TO36(-923), .W2TO37(-811), .W2TO38(-776), .W2TO39(379), .W2TO40(235), .W2TO41(148), .W2TO42(652), .W2TO43(490), .W2TO44(-546), .W2TO45(-823), .W2TO46(2), .W2TO47(-372), .W2TO48(-463), .W2TO49(19), .W2TO50(403), .W2TO51(814), .W2TO52(-91), .W2TO53(66), .W2TO54(618), .W2TO55(-221), .W2TO56(486), .W2TO57(970), .W2TO58(-578), .W2TO59(157), .W2TO60(441), .W2TO61(-732), .W2TO62(626), .W2TO63(474), .W3TO0(489), .W3TO1(687), .W3TO2(500), .W3TO3(482), .W3TO4(284), .W3TO5(279), .W3TO6(656), .W3TO7(668), .W3TO8(-556), .W3TO9(324), .W3TO10(-641), .W3TO11(643), .W3TO12(-935), .W3TO13(-931), .W3TO14(-960), .W3TO15(291), .W3TO16(63), .W3TO17(-944), .W3TO18(-946), .W3TO19(495), .W3TO20(497), .W3TO21(-536), .W3TO22(569), .W3TO23(688), .W3TO24(661), .W3TO25(110), .W3TO26(384), .W3TO27(544), .W3TO28(477), .W3TO29(-185), .W3TO30(343), .W3TO31(394), .W3TO32(630), .W3TO33(-300), .W3TO34(47), .W3TO35(-615), .W3TO36(-494), .W3TO37(83), .W3TO38(-396), .W3TO39(290), .W3TO40(-901), .W3TO41(-780), .W3TO42(515), .W3TO43(-113), .W3TO44(939), .W3TO45(-754), .W3TO46(-283), .W3TO47(847), .W3TO48(672), .W3TO49(956), .W3TO50(-608), .W3TO51(-280), .W3TO52(290), .W3TO53(-445), .W3TO54(-905), .W3TO55(163), .W3TO56(-624), .W3TO57(579), .W3TO58(-238), .W3TO59(-346), .W3TO60(303), .W3TO61(250), .W3TO62(-376), .W3TO63(496), .W4TO0(-193), .W4TO1(530), .W4TO2(-911), .W4TO3(820), .W4TO4(293), .W4TO5(-94), .W4TO6(-955), .W4TO7(-581), .W4TO8(227), .W4TO9(856), .W4TO10(208), .W4TO11(123), .W4TO12(-170), .W4TO13(672), .W4TO14(163), .W4TO15(489), .W4TO16(-507), .W4TO17(-770), .W4TO18(980), .W4TO19(-934), .W4TO20(-556), .W4TO21(-168), .W4TO22(-520), .W4TO23(-468), .W4TO24(112), .W4TO25(220), .W4TO26(214), .W4TO27(523), .W4TO28(-568), .W4TO29(787), .W4TO30(321), .W4TO31(-909), .W4TO32(194), .W4TO33(-244), .W4TO34(-310), .W4TO35(-601), .W4TO36(431), .W4TO37(955), .W4TO38(-443), .W4TO39(311), .W4TO40(-125), .W4TO41(-133), .W4TO42(-788), .W4TO43(-496), .W4TO44(736), .W4TO45(-767), .W4TO46(-366), .W4TO47(430), .W4TO48(-240), .W4TO49(-458), .W4TO50(894), .W4TO51(820), .W4TO52(221), .W4TO53(992), .W4TO54(973), .W4TO55(756), .W4TO56(3), .W4TO57(623), .W4TO58(592), .W4TO59(-644), .W4TO60(215), .W4TO61(-803), .W4TO62(-541), .W4TO63(-713), .W5TO0(-380), .W5TO1(-92), .W5TO2(-406), .W5TO3(119), .W5TO4(744), .W5TO5(-585), .W5TO6(-884), .W5TO7(816), .W5TO8(-319), .W5TO9(682), .W5TO10(865), .W5TO11(619), .W5TO12(-873), .W5TO13(-193), .W5TO14(-485), .W5TO15(288), .W5TO16(146), .W5TO17(851), .W5TO18(-211), .W5TO19(675), .W5TO20(364), .W5TO21(-332), .W5TO22(-431), .W5TO23(410), .W5TO24(143), .W5TO25(943), .W5TO26(-560), .W5TO27(-527), .W5TO28(387), .W5TO29(323), .W5TO30(840), .W5TO31(844), .W5TO32(-493), .W5TO33(75), .W5TO34(-208), .W5TO35(-816), .W5TO36(-453), .W5TO37(-827), .W5TO38(953), .W5TO39(800), .W5TO40(668), .W5TO41(959), .W5TO42(195), .W5TO43(360), .W5TO44(-556), .W5TO45(852), .W5TO46(-922), .W5TO47(264), .W5TO48(-920), .W5TO49(947), .W5TO50(751), .W5TO51(7), .W5TO52(179), .W5TO53(-437), .W5TO54(-693), .W5TO55(659), .W5TO56(-736), .W5TO57(-735), .W5TO58(-310), .W5TO59(976), .W5TO60(-32), .W5TO61(-384), .W5TO62(-499), .W5TO63(563), .W6TO0(-707), .W6TO1(-122), .W6TO2(736), .W6TO3(-971), .W6TO4(515), .W6TO5(958), .W6TO6(-533), .W6TO7(481), .W6TO8(601), .W6TO9(742), .W6TO10(392), .W6TO11(-557), .W6TO12(-836), .W6TO13(118), .W6TO14(119), .W6TO15(-200), .W6TO16(92), .W6TO17(-666), .W6TO18(-652), .W6TO19(430), .W6TO20(994), .W6TO21(602), .W6TO22(-667), .W6TO23(548), .W6TO24(-418), .W6TO25(855), .W6TO26(-53), .W6TO27(-203), .W6TO28(-800), .W6TO29(10), .W6TO30(-823), .W6TO31(369), .W6TO32(-724), .W6TO33(-59), .W6TO34(-504), .W6TO35(999), .W6TO36(-454), .W6TO37(170), .W6TO38(-970), .W6TO39(222), .W6TO40(22), .W6TO41(-33), .W6TO42(-193), .W6TO43(778), .W6TO44(-632), .W6TO45(387), .W6TO46(555), .W6TO47(469), .W6TO48(214), .W6TO49(401), .W6TO50(-518), .W6TO51(-829), .W6TO52(821), .W6TO53(71), .W6TO54(-516), .W6TO55(687), .W6TO56(632), .W6TO57(-522), .W6TO58(744), .W6TO59(-346), .W6TO60(-235), .W6TO61(-189), .W6TO62(12), .W6TO63(-518), .W7TO0(-51), .W7TO1(-475), .W7TO2(-217), .W7TO3(775), .W7TO4(-313), .W7TO5(-713), .W7TO6(451), .W7TO7(-424), .W7TO8(547), .W7TO9(994), .W7TO10(116), .W7TO11(-654), .W7TO12(-129), .W7TO13(-175), .W7TO14(-968), .W7TO15(-845), .W7TO16(376), .W7TO17(99), .W7TO18(865), .W7TO19(189), .W7TO20(380), .W7TO21(76), .W7TO22(156), .W7TO23(-922), .W7TO24(-489), .W7TO25(220), .W7TO26(-856), .W7TO27(-92), .W7TO28(484), .W7TO29(-942), .W7TO30(758), .W7TO31(480), .W7TO32(257), .W7TO33(-416), .W7TO34(-288), .W7TO35(-715), .W7TO36(-486), .W7TO37(348), .W7TO38(-945), .W7TO39(869), .W7TO40(-832), .W7TO41(-944), .W7TO42(-708), .W7TO43(753), .W7TO44(-615), .W7TO45(-457), .W7TO46(-115), .W7TO47(-869), .W7TO48(580), .W7TO49(-379), .W7TO50(591), .W7TO51(-235), .W7TO52(-858), .W7TO53(645), .W7TO54(343), .W7TO55(49), .W7TO56(-517), .W7TO57(893), .W7TO58(-36), .W7TO59(835), .W7TO60(589), .W7TO61(355), .W7TO62(34), .W7TO63(959), .W8TO0(-880), .W8TO1(741), .W8TO2(-904), .W8TO3(-206), .W8TO4(143), .W8TO5(-28), .W8TO6(-142), .W8TO7(-123), .W8TO8(-776), .W8TO9(-720), .W8TO10(-395), .W8TO11(784), .W8TO12(561), .W8TO13(-567), .W8TO14(-814), .W8TO15(38), .W8TO16(-643), .W8TO17(-382), .W8TO18(-663), .W8TO19(-305), .W8TO20(220), .W8TO21(950), .W8TO22(333), .W8TO23(-183), .W8TO24(-302), .W8TO25(-275), .W8TO26(802), .W8TO27(-319), .W8TO28(-872), .W8TO29(2), .W8TO30(-826), .W8TO31(-835), .W8TO32(925), .W8TO33(-83), .W8TO34(881), .W8TO35(477), .W8TO36(281), .W8TO37(-80), .W8TO38(-842), .W8TO39(428), .W8TO40(-396), .W8TO41(549), .W8TO42(-385), .W8TO43(-12), .W8TO44(261), .W8TO45(-657), .W8TO46(255), .W8TO47(-775), .W8TO48(-290), .W8TO49(-196), .W8TO50(-523), .W8TO51(966), .W8TO52(-876), .W8TO53(778), .W8TO54(269), .W8TO55(921), .W8TO56(164), .W8TO57(421), .W8TO58(712), .W8TO59(605), .W8TO60(-607), .W8TO61(38), .W8TO62(-329), .W8TO63(879), .W9TO0(290), .W9TO1(38), .W9TO2(326), .W9TO3(-746), .W9TO4(699), .W9TO5(-377), .W9TO6(-830), .W9TO7(-440), .W9TO8(253), .W9TO9(-474), .W9TO10(-852), .W9TO11(934), .W9TO12(349), .W9TO13(-696), .W9TO14(293), .W9TO15(-768), .W9TO16(-670), .W9TO17(-763), .W9TO18(-176), .W9TO19(946), .W9TO20(-728), .W9TO21(-743), .W9TO22(-665), .W9TO23(268), .W9TO24(376), .W9TO25(236), .W9TO26(-946), .W9TO27(176), .W9TO28(-910), .W9TO29(274), .W9TO30(-314), .W9TO31(923), .W9TO32(753), .W9TO33(510), .W9TO34(658), .W9TO35(50), .W9TO36(-191), .W9TO37(-785), .W9TO38(-3), .W9TO39(-636), .W9TO40(568), .W9TO41(-703), .W9TO42(-754), .W9TO43(692), .W9TO44(878), .W9TO45(-100), .W9TO46(-701), .W9TO47(97), .W9TO48(-695), .W9TO49(-387), .W9TO50(866), .W9TO51(-862), .W9TO52(-901), .W9TO53(-778), .W9TO54(-74), .W9TO55(-583), .W9TO56(815), .W9TO57(-290), .W9TO58(-219), .W9TO59(-384), .W9TO60(166), .W9TO61(749), .W9TO62(-698), .W9TO63(431), .W10TO0(528), .W10TO1(476), .W10TO2(-675), .W10TO3(132), .W10TO4(183), .W10TO5(-896), .W10TO6(-21), .W10TO7(501), .W10TO8(-913), .W10TO9(177), .W10TO10(210), .W10TO11(-577), .W10TO12(-852), .W10TO13(292), .W10TO14(569), .W10TO15(151), .W10TO16(-517), .W10TO17(-638), .W10TO18(-714), .W10TO19(1), .W10TO20(-771), .W10TO21(-874), .W10TO22(-756), .W10TO23(-822), .W10TO24(322), .W10TO25(-182), .W10TO26(294), .W10TO27(-277), .W10TO28(428), .W10TO29(-5), .W10TO30(582), .W10TO31(917), .W10TO32(-542), .W10TO33(-549), .W10TO34(74), .W10TO35(-353), .W10TO36(532), .W10TO37(637), .W10TO38(-68), .W10TO39(-904), .W10TO40(759), .W10TO41(779), .W10TO42(892), .W10TO43(622), .W10TO44(798), .W10TO45(900), .W10TO46(755), .W10TO47(920), .W10TO48(-105), .W10TO49(680), .W10TO50(-493), .W10TO51(551), .W10TO52(848), .W10TO53(-293), .W10TO54(-381), .W10TO55(467), .W10TO56(541), .W10TO57(-65), .W10TO58(231), .W10TO59(349), .W10TO60(-981), .W10TO61(-261), .W10TO62(-487), .W10TO63(686), .W11TO0(-558), .W11TO1(963), .W11TO2(992), .W11TO3(207), .W11TO4(-627), .W11TO5(66), .W11TO6(980), .W11TO7(-282), .W11TO8(-650), .W11TO9(718), .W11TO10(623), .W11TO11(-997), .W11TO12(-228), .W11TO13(563), .W11TO14(-83), .W11TO15(378), .W11TO16(714), .W11TO17(245), .W11TO18(529), .W11TO19(266), .W11TO20(-924), .W11TO21(-515), .W11TO22(404), .W11TO23(-801), .W11TO24(592), .W11TO25(-647), .W11TO26(-971), .W11TO27(27), .W11TO28(56), .W11TO29(-39), .W11TO30(-500), .W11TO31(-736), .W11TO32(-121), .W11TO33(-670), .W11TO34(-985), .W11TO35(830), .W11TO36(-169), .W11TO37(814), .W11TO38(147), .W11TO39(-278), .W11TO40(230), .W11TO41(754), .W11TO42(-643), .W11TO43(-505), .W11TO44(-51), .W11TO45(-553), .W11TO46(-6), .W11TO47(-175), .W11TO48(-328), .W11TO49(-226), .W11TO50(990), .W11TO51(-4), .W11TO52(-910), .W11TO53(997), .W11TO54(625), .W11TO55(-352), .W11TO56(-153), .W11TO57(477), .W11TO58(-310), .W11TO59(-151), .W11TO60(-299), .W11TO61(-79), .W11TO62(62), .W11TO63(896), .W12TO0(-432), .W12TO1(499), .W12TO2(-681), .W12TO3(-736), .W12TO4(-150), .W12TO5(666), .W12TO6(-363), .W12TO7(734), .W12TO8(-597), .W12TO9(-332), .W12TO10(170), .W12TO11(488), .W12TO12(345), .W12TO13(-490), .W12TO14(455), .W12TO15(-410), .W12TO16(-545), .W12TO17(-801), .W12TO18(-291), .W12TO19(742), .W12TO20(588), .W12TO21(-632), .W12TO22(-468), .W12TO23(402), .W12TO24(963), .W12TO25(184), .W12TO26(-420), .W12TO27(-938), .W12TO28(-57), .W12TO29(-858), .W12TO30(-710), .W12TO31(666), .W12TO32(759), .W12TO33(376), .W12TO34(-974), .W12TO35(-352), .W12TO36(832), .W12TO37(974), .W12TO38(313), .W12TO39(593), .W12TO40(119), .W12TO41(-88), .W12TO42(-197), .W12TO43(274), .W12TO44(-896), .W12TO45(198), .W12TO46(557), .W12TO47(-695), .W12TO48(-315), .W12TO49(-834), .W12TO50(-864), .W12TO51(-533), .W12TO52(-945), .W12TO53(636), .W12TO54(354), .W12TO55(324), .W12TO56(934), .W12TO57(-56), .W12TO58(314), .W12TO59(532), .W12TO60(-741), .W12TO61(374), .W12TO62(468), .W12TO63(80), .W13TO0(813), .W13TO1(-41), .W13TO2(700), .W13TO3(689), .W13TO4(699), .W13TO5(824), .W13TO6(460), .W13TO7(691), .W13TO8(-253), .W13TO9(-114), .W13TO10(502), .W13TO11(-391), .W13TO12(-207), .W13TO13(-575), .W13TO14(-170), .W13TO15(-418), .W13TO16(110), .W13TO17(-196), .W13TO18(-741), .W13TO19(-968), .W13TO20(727), .W13TO21(-500), .W13TO22(-106), .W13TO23(-369), .W13TO24(-777), .W13TO25(934), .W13TO26(-27), .W13TO27(570), .W13TO28(-414), .W13TO29(-413), .W13TO30(-693), .W13TO31(-399), .W13TO32(-710), .W13TO33(940), .W13TO34(703), .W13TO35(-250), .W13TO36(614), .W13TO37(774), .W13TO38(-993), .W13TO39(1), .W13TO40(-897), .W13TO41(-96), .W13TO42(621), .W13TO43(418), .W13TO44(364), .W13TO45(387), .W13TO46(606), .W13TO47(497), .W13TO48(-58), .W13TO49(534), .W13TO50(-326), .W13TO51(-771), .W13TO52(45), .W13TO53(454), .W13TO54(688), .W13TO55(-989), .W13TO56(-957), .W13TO57(-142), .W13TO58(-535), .W13TO59(-288), .W13TO60(-812), .W13TO61(448), .W13TO62(-767), .W13TO63(41), .W14TO0(939), .W14TO1(720), .W14TO2(-820), .W14TO3(-865), .W14TO4(155), .W14TO5(-22), .W14TO6(-416), .W14TO7(-225), .W14TO8(827), .W14TO9(-616), .W14TO10(744), .W14TO11(882), .W14TO12(811), .W14TO13(-271), .W14TO14(-288), .W14TO15(855), .W14TO16(840), .W14TO17(-317), .W14TO18(-680), .W14TO19(358), .W14TO20(-129), .W14TO21(66), .W14TO22(310), .W14TO23(896), .W14TO24(-47), .W14TO25(-148), .W14TO26(-493), .W14TO27(-68), .W14TO28(132), .W14TO29(28), .W14TO30(-734), .W14TO31(760), .W14TO32(-340), .W14TO33(-996), .W14TO34(-200), .W14TO35(-851), .W14TO36(-916), .W14TO37(-166), .W14TO38(497), .W14TO39(604), .W14TO40(246), .W14TO41(-606), .W14TO42(-282), .W14TO43(194), .W14TO44(914), .W14TO45(651), .W14TO46(842), .W14TO47(-40), .W14TO48(-653), .W14TO49(-994), .W14TO50(-205), .W14TO51(113), .W14TO52(651), .W14TO53(-962), .W14TO54(573), .W14TO55(-331), .W14TO56(402), .W14TO57(161), .W14TO58(996), .W14TO59(-306), .W14TO60(543), .W14TO61(-569), .W14TO62(598), .W14TO63(-22), .W15TO0(-467), .W15TO1(-837), .W15TO2(800), .W15TO3(574), .W15TO4(773), .W15TO5(-573), .W15TO6(0), .W15TO7(-880), .W15TO8(-735), .W15TO9(839), .W15TO10(230), .W15TO11(46), .W15TO12(-510), .W15TO13(280), .W15TO14(-846), .W15TO15(-132), .W15TO16(-557), .W15TO17(265), .W15TO18(108), .W15TO19(965), .W15TO20(69), .W15TO21(635), .W15TO22(691), .W15TO23(692), .W15TO24(183), .W15TO25(649), .W15TO26(432), .W15TO27(284), .W15TO28(435), .W15TO29(-537), .W15TO30(970), .W15TO31(-519), .W15TO32(507), .W15TO33(691), .W15TO34(186), .W15TO35(308), .W15TO36(432), .W15TO37(140), .W15TO38(671), .W15TO39(965), .W15TO40(472), .W15TO41(-185), .W15TO42(245), .W15TO43(-927), .W15TO44(112), .W15TO45(-29), .W15TO46(-861), .W15TO47(-524), .W15TO48(-365), .W15TO49(589), .W15TO50(-948), .W15TO51(890), .W15TO52(368), .W15TO53(-421), .W15TO54(-738), .W15TO55(189), .W15TO56(483), .W15TO57(169), .W15TO58(-790), .W15TO59(971), .W15TO60(76), .W15TO61(-437), .W15TO62(234), .W15TO63(-873), .W16TO0(-934), .W16TO1(608), .W16TO2(-475), .W16TO3(896), .W16TO4(-869), .W16TO5(-74), .W16TO6(-480), .W16TO7(275), .W16TO8(161), .W16TO9(-216), .W16TO10(48), .W16TO11(-692), .W16TO12(-522), .W16TO13(731), .W16TO14(723), .W16TO15(974), .W16TO16(-123), .W16TO17(-868), .W16TO18(-349), .W16TO19(-827), .W16TO20(563), .W16TO21(651), .W16TO22(-938), .W16TO23(329), .W16TO24(404), .W16TO25(-521), .W16TO26(-120), .W16TO27(997), .W16TO28(751), .W16TO29(353), .W16TO30(271), .W16TO31(689), .W16TO32(-264), .W16TO33(-179), .W16TO34(891), .W16TO35(-81), .W16TO36(-325), .W16TO37(345), .W16TO38(-118), .W16TO39(506), .W16TO40(-217), .W16TO41(211), .W16TO42(-619), .W16TO43(-736), .W16TO44(768), .W16TO45(985), .W16TO46(-498), .W16TO47(-371), .W16TO48(-396), .W16TO49(366), .W16TO50(-670), .W16TO51(437), .W16TO52(203), .W16TO53(-796), .W16TO54(201), .W16TO55(537), .W16TO56(-879), .W16TO57(-862), .W16TO58(994), .W16TO59(345), .W16TO60(-927), .W16TO61(-107), .W16TO62(90), .W16TO63(-158), .W17TO0(251), .W17TO1(642), .W17TO2(-209), .W17TO3(-499), .W17TO4(36), .W17TO5(-986), .W17TO6(-589), .W17TO7(320), .W17TO8(-425), .W17TO9(-446), .W17TO10(145), .W17TO11(-131), .W17TO12(-711), .W17TO13(990), .W17TO14(937), .W17TO15(-56), .W17TO16(480), .W17TO17(324), .W17TO18(431), .W17TO19(34), .W17TO20(-505), .W17TO21(7), .W17TO22(911), .W17TO23(423), .W17TO24(-983), .W17TO25(-181), .W17TO26(-129), .W17TO27(754), .W17TO28(-142), .W17TO29(-355), .W17TO30(542), .W17TO31(839), .W17TO32(-695), .W17TO33(995), .W17TO34(846), .W17TO35(-335), .W17TO36(19), .W17TO37(-743), .W17TO38(840), .W17TO39(-151), .W17TO40(-539), .W17TO41(-579), .W17TO42(150), .W17TO43(756), .W17TO44(-245), .W17TO45(262), .W17TO46(697), .W17TO47(-953), .W17TO48(594), .W17TO49(701), .W17TO50(-476), .W17TO51(-560), .W17TO52(161), .W17TO53(172), .W17TO54(-598), .W17TO55(-67), .W17TO56(108), .W17TO57(-635), .W17TO58(-351), .W17TO59(213), .W17TO60(-652), .W17TO61(-114), .W17TO62(-108), .W17TO63(839), .W18TO0(444), .W18TO1(366), .W18TO2(-489), .W18TO3(364), .W18TO4(-981), .W18TO5(-156), .W18TO6(955), .W18TO7(-343), .W18TO8(869), .W18TO9(540), .W18TO10(-442), .W18TO11(-519), .W18TO12(-696), .W18TO13(47), .W18TO14(46), .W18TO15(-183), .W18TO16(646), .W18TO17(656), .W18TO18(63), .W18TO19(381), .W18TO20(-13), .W18TO21(-39), .W18TO22(233), .W18TO23(-565), .W18TO24(-738), .W18TO25(124), .W18TO26(-377), .W18TO27(-18), .W18TO28(-415), .W18TO29(-469), .W18TO30(-154), .W18TO31(-995), .W18TO32(-458), .W18TO33(-262), .W18TO34(-17), .W18TO35(892), .W18TO36(112), .W18TO37(720), .W18TO38(195), .W18TO39(-185), .W18TO40(-964), .W18TO41(859), .W18TO42(-279), .W18TO43(806), .W18TO44(655), .W18TO45(-854), .W18TO46(-738), .W18TO47(-433), .W18TO48(-81), .W18TO49(286), .W18TO50(778), .W18TO51(-141), .W18TO52(487), .W18TO53(827), .W18TO54(-733), .W18TO55(886), .W18TO56(593), .W18TO57(491), .W18TO58(-107), .W18TO59(-851), .W18TO60(-479), .W18TO61(320), .W18TO62(-951), .W18TO63(543), .W19TO0(946), .W19TO1(-753), .W19TO2(290), .W19TO3(698), .W19TO4(408), .W19TO5(691), .W19TO6(865), .W19TO7(617), .W19TO8(-97), .W19TO9(167), .W19TO10(-24), .W19TO11(227), .W19TO12(29), .W19TO13(280), .W19TO14(595), .W19TO15(910), .W19TO16(5), .W19TO17(-101), .W19TO18(-527), .W19TO19(801), .W19TO20(603), .W19TO21(-243), .W19TO22(-624), .W19TO23(-109), .W19TO24(880), .W19TO25(-247), .W19TO26(-359), .W19TO27(776), .W19TO28(793), .W19TO29(-250), .W19TO30(899), .W19TO31(676), .W19TO32(175), .W19TO33(-508), .W19TO34(-526), .W19TO35(-340), .W19TO36(962), .W19TO37(121), .W19TO38(540), .W19TO39(-100), .W19TO40(732), .W19TO41(907), .W19TO42(390), .W19TO43(40), .W19TO44(-622), .W19TO45(630), .W19TO46(688), .W19TO47(888), .W19TO48(728), .W19TO49(-184), .W19TO50(-396), .W19TO51(-51), .W19TO52(953), .W19TO53(662), .W19TO54(-743), .W19TO55(673), .W19TO56(-209), .W19TO57(953), .W19TO58(999), .W19TO59(463), .W19TO60(679), .W19TO61(-572), .W19TO62(-288), .W19TO63(690), .W20TO0(-362), .W20TO1(-10), .W20TO2(530), .W20TO3(-116), .W20TO4(145), .W20TO5(126), .W20TO6(758), .W20TO7(583), .W20TO8(516), .W20TO9(-343), .W20TO10(-56), .W20TO11(909), .W20TO12(-719), .W20TO13(378), .W20TO14(-614), .W20TO15(-473), .W20TO16(-153), .W20TO17(-495), .W20TO18(-29), .W20TO19(426), .W20TO20(-219), .W20TO21(-763), .W20TO22(225), .W20TO23(870), .W20TO24(460), .W20TO25(298), .W20TO26(-778), .W20TO27(161), .W20TO28(-476), .W20TO29(-211), .W20TO30(-10), .W20TO31(-390), .W20TO32(954), .W20TO33(-745), .W20TO34(252), .W20TO35(955), .W20TO36(-157), .W20TO37(38), .W20TO38(-697), .W20TO39(970), .W20TO40(585), .W20TO41(247), .W20TO42(366), .W20TO43(-933), .W20TO44(282), .W20TO45(359), .W20TO46(720), .W20TO47(288), .W20TO48(8), .W20TO49(777), .W20TO50(531), .W20TO51(-489), .W20TO52(495), .W20TO53(488), .W20TO54(145), .W20TO55(146), .W20TO56(-173), .W20TO57(810), .W20TO58(740), .W20TO59(360), .W20TO60(869), .W20TO61(659), .W20TO62(81), .W20TO63(-494), .W21TO0(130), .W21TO1(292), .W21TO2(621), .W21TO3(66), .W21TO4(948), .W21TO5(-583), .W21TO6(-534), .W21TO7(266), .W21TO8(203), .W21TO9(-377), .W21TO10(273), .W21TO11(943), .W21TO12(829), .W21TO13(601), .W21TO14(-587), .W21TO15(738), .W21TO16(159), .W21TO17(505), .W21TO18(28), .W21TO19(-832), .W21TO20(-799), .W21TO21(427), .W21TO22(275), .W21TO23(-510), .W21TO24(-851), .W21TO25(-743), .W21TO26(553), .W21TO27(-930), .W21TO28(290), .W21TO29(846), .W21TO30(-782), .W21TO31(884), .W21TO32(357), .W21TO33(-281), .W21TO34(-614), .W21TO35(226), .W21TO36(13), .W21TO37(-231), .W21TO38(20), .W21TO39(-7), .W21TO40(866), .W21TO41(-446), .W21TO42(685), .W21TO43(873), .W21TO44(524), .W21TO45(890), .W21TO46(-659), .W21TO47(-965), .W21TO48(-9), .W21TO49(-586), .W21TO50(-393), .W21TO51(532), .W21TO52(-159), .W21TO53(439), .W21TO54(361), .W21TO55(712), .W21TO56(-231), .W21TO57(877), .W21TO58(922), .W21TO59(23), .W21TO60(-509), .W21TO61(-619), .W21TO62(18), .W21TO63(-440), .W22TO0(-781), .W22TO1(-885), .W22TO2(363), .W22TO3(122), .W22TO4(95), .W22TO5(-732), .W22TO6(688), .W22TO7(-723), .W22TO8(-372), .W22TO9(474), .W22TO10(-106), .W22TO11(838), .W22TO12(514), .W22TO13(429), .W22TO14(-544), .W22TO15(-473), .W22TO16(-298), .W22TO17(839), .W22TO18(312), .W22TO19(700), .W22TO20(-62), .W22TO21(-778), .W22TO22(-375), .W22TO23(440), .W22TO24(-655), .W22TO25(-850), .W22TO26(-993), .W22TO27(-706), .W22TO28(285), .W22TO29(36), .W22TO30(-212), .W22TO31(-798), .W22TO32(-573), .W22TO33(811), .W22TO34(-615), .W22TO35(105), .W22TO36(-203), .W22TO37(-613), .W22TO38(619), .W22TO39(-612), .W22TO40(863), .W22TO41(-240), .W22TO42(435), .W22TO43(-823), .W22TO44(-883), .W22TO45(-586), .W22TO46(-30), .W22TO47(886), .W22TO48(-711), .W22TO49(991), .W22TO50(-43), .W22TO51(331), .W22TO52(7), .W22TO53(130), .W22TO54(466), .W22TO55(-459), .W22TO56(563), .W22TO57(-480), .W22TO58(543), .W22TO59(397), .W22TO60(-20), .W22TO61(849), .W22TO62(-747), .W22TO63(-975), .W23TO0(693), .W23TO1(-844), .W23TO2(887), .W23TO3(-847), .W23TO4(-388), .W23TO5(-638), .W23TO6(-751), .W23TO7(-593), .W23TO8(436), .W23TO9(310), .W23TO10(26), .W23TO11(-154), .W23TO12(520), .W23TO13(-24), .W23TO14(832), .W23TO15(545), .W23TO16(424), .W23TO17(-766), .W23TO18(-313), .W23TO19(-249), .W23TO20(-74), .W23TO21(-407), .W23TO22(-433), .W23TO23(938), .W23TO24(-209), .W23TO25(405), .W23TO26(920), .W23TO27(-181), .W23TO28(328), .W23TO29(684), .W23TO30(-496), .W23TO31(-578), .W23TO32(-853), .W23TO33(107), .W23TO34(408), .W23TO35(505), .W23TO36(270), .W23TO37(-873), .W23TO38(-975), .W23TO39(-552), .W23TO40(-394), .W23TO41(67), .W23TO42(114), .W23TO43(-356), .W23TO44(331), .W23TO45(-628), .W23TO46(233), .W23TO47(-290), .W23TO48(-394), .W23TO49(-518), .W23TO50(331), .W23TO51(-672), .W23TO52(-860), .W23TO53(-658), .W23TO54(865), .W23TO55(338), .W23TO56(192), .W23TO57(416), .W23TO58(325), .W23TO59(737), .W23TO60(832), .W23TO61(653), .W23TO62(155), .W23TO63(61), .W24TO0(-706), .W24TO1(205), .W24TO2(-213), .W24TO3(-902), .W24TO4(520), .W24TO5(334), .W24TO6(-84), .W24TO7(351), .W24TO8(-149), .W24TO9(536), .W24TO10(852), .W24TO11(-360), .W24TO12(-406), .W24TO13(-92), .W24TO14(-566), .W24TO15(-558), .W24TO16(185), .W24TO17(-404), .W24TO18(-123), .W24TO19(676), .W24TO20(378), .W24TO21(638), .W24TO22(-590), .W24TO23(716), .W24TO24(84), .W24TO25(853), .W24TO26(-410), .W24TO27(831), .W24TO28(-842), .W24TO29(-464), .W24TO30(709), .W24TO31(228), .W24TO32(-38), .W24TO33(376), .W24TO34(-58), .W24TO35(428), .W24TO36(-103), .W24TO37(-701), .W24TO38(109), .W24TO39(-219), .W24TO40(249), .W24TO41(961), .W24TO42(-762), .W24TO43(-63), .W24TO44(-737), .W24TO45(-62), .W24TO46(-555), .W24TO47(-214), .W24TO48(760), .W24TO49(-373), .W24TO50(-572), .W24TO51(758), .W24TO52(-407), .W24TO53(-748), .W24TO54(-52), .W24TO55(447), .W24TO56(507), .W24TO57(640), .W24TO58(-996), .W24TO59(-816), .W24TO60(-984), .W24TO61(498), .W24TO62(719), .W24TO63(-122), .W25TO0(-945), .W25TO1(829), .W25TO2(-173), .W25TO3(-169), .W25TO4(386), .W25TO5(874), .W25TO6(232), .W25TO7(383), .W25TO8(471), .W25TO9(-5), .W25TO10(-280), .W25TO11(-231), .W25TO12(676), .W25TO13(-793), .W25TO14(664), .W25TO15(-330), .W25TO16(-286), .W25TO17(-239), .W25TO18(662), .W25TO19(434), .W25TO20(-805), .W25TO21(-308), .W25TO22(-925), .W25TO23(565), .W25TO24(-4), .W25TO25(379), .W25TO26(-847), .W25TO27(820), .W25TO28(269), .W25TO29(781), .W25TO30(-665), .W25TO31(-328), .W25TO32(-549), .W25TO33(49), .W25TO34(425), .W25TO35(-310), .W25TO36(749), .W25TO37(-948), .W25TO38(-412), .W25TO39(4), .W25TO40(377), .W25TO41(-376), .W25TO42(893), .W25TO43(-511), .W25TO44(-309), .W25TO45(-310), .W25TO46(-325), .W25TO47(-884), .W25TO48(-527), .W25TO49(-148), .W25TO50(-522), .W25TO51(-423), .W25TO52(565), .W25TO53(322), .W25TO54(52), .W25TO55(319), .W25TO56(838), .W25TO57(741), .W25TO58(853), .W25TO59(-797), .W25TO60(436), .W25TO61(540), .W25TO62(915), .W25TO63(-947), .W26TO0(-225), .W26TO1(-535), .W26TO2(-750), .W26TO3(-818), .W26TO4(69), .W26TO5(724), .W26TO6(-531), .W26TO7(-174), .W26TO8(-546), .W26TO9(-122), .W26TO10(391), .W26TO11(396), .W26TO12(411), .W26TO13(-274), .W26TO14(-882), .W26TO15(244), .W26TO16(-195), .W26TO17(324), .W26TO18(-468), .W26TO19(913), .W26TO20(-495), .W26TO21(125), .W26TO22(211), .W26TO23(-144), .W26TO24(632), .W26TO25(102), .W26TO26(30), .W26TO27(-777), .W26TO28(-447), .W26TO29(599), .W26TO30(714), .W26TO31(-566), .W26TO32(997), .W26TO33(-903), .W26TO34(-243), .W26TO35(-864), .W26TO36(-229), .W26TO37(987), .W26TO38(-810), .W26TO39(-749), .W26TO40(829), .W26TO41(-293), .W26TO42(-319), .W26TO43(-145), .W26TO44(328), .W26TO45(144), .W26TO46(-443), .W26TO47(478), .W26TO48(-395), .W26TO49(722), .W26TO50(233), .W26TO51(-958), .W26TO52(-462), .W26TO53(-603), .W26TO54(-280), .W26TO55(284), .W26TO56(-354), .W26TO57(-856), .W26TO58(836), .W26TO59(-827), .W26TO60(-827), .W26TO61(667), .W26TO62(-976), .W26TO63(994), .W27TO0(679), .W27TO1(-405), .W27TO2(-295), .W27TO3(864), .W27TO4(-753), .W27TO5(106), .W27TO6(586), .W27TO7(-746), .W27TO8(-107), .W27TO9(-86), .W27TO10(914), .W27TO11(41), .W27TO12(985), .W27TO13(-885), .W27TO14(-451), .W27TO15(-430), .W27TO16(465), .W27TO17(-887), .W27TO18(518), .W27TO19(633), .W27TO20(-65), .W27TO21(-521), .W27TO22(-386), .W27TO23(411), .W27TO24(-80), .W27TO25(-551), .W27TO26(445), .W27TO27(607), .W27TO28(825), .W27TO29(199), .W27TO30(479), .W27TO31(-886), .W27TO32(404), .W27TO33(-278), .W27TO34(-993), .W27TO35(528), .W27TO36(775), .W27TO37(-513), .W27TO38(-775), .W27TO39(659), .W27TO40(191), .W27TO41(-448), .W27TO42(832), .W27TO43(-990), .W27TO44(-157), .W27TO45(-465), .W27TO46(521), .W27TO47(-745), .W27TO48(461), .W27TO49(-563), .W27TO50(-996), .W27TO51(427), .W27TO52(-101), .W27TO53(860), .W27TO54(-668), .W27TO55(147), .W27TO56(200), .W27TO57(-323), .W27TO58(429), .W27TO59(346), .W27TO60(730), .W27TO61(-933), .W27TO62(268), .W27TO63(584), .W28TO0(934), .W28TO1(-930), .W28TO2(-207), .W28TO3(340), .W28TO4(696), .W28TO5(-388), .W28TO6(-361), .W28TO7(569), .W28TO8(-766), .W28TO9(231), .W28TO10(761), .W28TO11(-101), .W28TO12(74), .W28TO13(130), .W28TO14(-690), .W28TO15(552), .W28TO16(417), .W28TO17(614), .W28TO18(688), .W28TO19(172), .W28TO20(-692), .W28TO21(415), .W28TO22(-926), .W28TO23(365), .W28TO24(-496), .W28TO25(-81), .W28TO26(-273), .W28TO27(-897), .W28TO28(681), .W28TO29(477), .W28TO30(-203), .W28TO31(565), .W28TO32(81), .W28TO33(866), .W28TO34(668), .W28TO35(-755), .W28TO36(-34), .W28TO37(-199), .W28TO38(731), .W28TO39(880), .W28TO40(-546), .W28TO41(-74), .W28TO42(-813), .W28TO43(390), .W28TO44(627), .W28TO45(-717), .W28TO46(-702), .W28TO47(207), .W28TO48(870), .W28TO49(-222), .W28TO50(-427), .W28TO51(-188), .W28TO52(831), .W28TO53(340), .W28TO54(-405), .W28TO55(209), .W28TO56(357), .W28TO57(-297), .W28TO58(530), .W28TO59(895), .W28TO60(-631), .W28TO61(-501), .W28TO62(172), .W28TO63(-435), .W29TO0(792), .W29TO1(523), .W29TO2(-447), .W29TO3(875), .W29TO4(292), .W29TO5(634), .W29TO6(-53), .W29TO7(597), .W29TO8(-368), .W29TO9(466), .W29TO10(-11), .W29TO11(-647), .W29TO12(-957), .W29TO13(-964), .W29TO14(868), .W29TO15(204), .W29TO16(579), .W29TO17(518), .W29TO18(-687), .W29TO19(-12), .W29TO20(684), .W29TO21(-878), .W29TO22(-792), .W29TO23(329), .W29TO24(744), .W29TO25(-842), .W29TO26(722), .W29TO27(199), .W29TO28(752), .W29TO29(-404), .W29TO30(-390), .W29TO31(925), .W29TO32(-394), .W29TO33(-310), .W29TO34(-435), .W29TO35(-895), .W29TO36(468), .W29TO37(-135), .W29TO38(546), .W29TO39(474), .W29TO40(462), .W29TO41(604), .W29TO42(-733), .W29TO43(28), .W29TO44(280), .W29TO45(787), .W29TO46(611), .W29TO47(-435), .W29TO48(-553), .W29TO49(806), .W29TO50(-401), .W29TO51(-493), .W29TO52(-888), .W29TO53(993), .W29TO54(618), .W29TO55(568), .W29TO56(-937), .W29TO57(63), .W29TO58(67), .W29TO59(566), .W29TO60(689), .W29TO61(704), .W29TO62(-54), .W29TO63(590), .W30TO0(949), .W30TO1(-878), .W30TO2(739), .W30TO3(-262), .W30TO4(-139), .W30TO5(-983), .W30TO6(310), .W30TO7(173), .W30TO8(980), .W30TO9(478), .W30TO10(28), .W30TO11(0), .W30TO12(502), .W30TO13(-811), .W30TO14(928), .W30TO15(-663), .W30TO16(-407), .W30TO17(-744), .W30TO18(112), .W30TO19(-632), .W30TO20(-515), .W30TO21(-963), .W30TO22(-664), .W30TO23(-163), .W30TO24(22), .W30TO25(-505), .W30TO26(239), .W30TO27(-396), .W30TO28(474), .W30TO29(-69), .W30TO30(739), .W30TO31(604), .W30TO32(-472), .W30TO33(331), .W30TO34(-231), .W30TO35(-405), .W30TO36(597), .W30TO37(400), .W30TO38(-794), .W30TO39(-947), .W30TO40(-534), .W30TO41(938), .W30TO42(528), .W30TO43(551), .W30TO44(-963), .W30TO45(-540), .W30TO46(-593), .W30TO47(691), .W30TO48(859), .W30TO49(-814), .W30TO50(-17), .W30TO51(491), .W30TO52(458), .W30TO53(346), .W30TO54(-226), .W30TO55(432), .W30TO56(764), .W30TO57(65), .W30TO58(-427), .W30TO59(724), .W30TO60(789), .W30TO61(-329), .W30TO62(979), .W30TO63(188), .W31TO0(837), .W31TO1(-152), .W31TO2(243), .W31TO3(-395), .W31TO4(178), .W31TO5(-591), .W31TO6(-592), .W31TO7(425), .W31TO8(-35), .W31TO9(-131), .W31TO10(-611), .W31TO11(930), .W31TO12(474), .W31TO13(-449), .W31TO14(-61), .W31TO15(-637), .W31TO16(799), .W31TO17(482), .W31TO18(327), .W31TO19(-947), .W31TO20(-58), .W31TO21(-926), .W31TO22(-993), .W31TO23(633), .W31TO24(-553), .W31TO25(-230), .W31TO26(-819), .W31TO27(65), .W31TO28(760), .W31TO29(-162), .W31TO30(762), .W31TO31(-81), .W31TO32(905), .W31TO33(-390), .W31TO34(-739), .W31TO35(98), .W31TO36(-533), .W31TO37(-488), .W31TO38(3), .W31TO39(-922), .W31TO40(-601), .W31TO41(-70), .W31TO42(461), .W31TO43(-223), .W31TO44(470), .W31TO45(-993), .W31TO46(-191), .W31TO47(-511), .W31TO48(-925), .W31TO49(-895), .W31TO50(-254), .W31TO51(-142), .W31TO52(285), .W31TO53(659), .W31TO54(-687), .W31TO55(497), .W31TO56(-561), .W31TO57(-781), .W31TO58(894), .W31TO59(476), .W31TO60(58), .W31TO61(611), .W31TO62(309), .W31TO63(87), .W32TO0(-428), .W32TO1(-138), .W32TO2(589), .W32TO3(-943), .W32TO4(443), .W32TO5(423), .W32TO6(169), .W32TO7(490), .W32TO8(297), .W32TO9(688), .W32TO10(-297), .W32TO11(332), .W32TO12(419), .W32TO13(-743), .W32TO14(-747), .W32TO15(840), .W32TO16(-573), .W32TO17(-356), .W32TO18(-691), .W32TO19(-324), .W32TO20(568), .W32TO21(400), .W32TO22(422), .W32TO23(696), .W32TO24(974), .W32TO25(-272), .W32TO26(-387), .W32TO27(-167), .W32TO28(-26), .W32TO29(969), .W32TO30(529), .W32TO31(162), .W32TO32(-719), .W32TO33(816), .W32TO34(-575), .W32TO35(857), .W32TO36(-357), .W32TO37(-363), .W32TO38(-28), .W32TO39(-524), .W32TO40(728), .W32TO41(767), .W32TO42(653), .W32TO43(-447), .W32TO44(82), .W32TO45(740), .W32TO46(-598), .W32TO47(-496), .W32TO48(-875), .W32TO49(-822), .W32TO50(-385), .W32TO51(-153), .W32TO52(673), .W32TO53(395), .W32TO54(867), .W32TO55(531), .W32TO56(341), .W32TO57(-589), .W32TO58(-517), .W32TO59(110), .W32TO60(612), .W32TO61(-547), .W32TO62(-460), .W32TO63(331), .W33TO0(158), .W33TO1(418), .W33TO2(687), .W33TO3(-752), .W33TO4(-543), .W33TO5(-285), .W33TO6(-787), .W33TO7(-483), .W33TO8(-790), .W33TO9(-536), .W33TO10(467), .W33TO11(-329), .W33TO12(28), .W33TO13(368), .W33TO14(666), .W33TO15(-851), .W33TO16(251), .W33TO17(-625), .W33TO18(824), .W33TO19(-188), .W33TO20(-20), .W33TO21(-110), .W33TO22(650), .W33TO23(533), .W33TO24(200), .W33TO25(770), .W33TO26(-546), .W33TO27(176), .W33TO28(87), .W33TO29(-859), .W33TO30(70), .W33TO31(-897), .W33TO32(-151), .W33TO33(-556), .W33TO34(524), .W33TO35(59), .W33TO36(-96), .W33TO37(138), .W33TO38(-848), .W33TO39(507), .W33TO40(733), .W33TO41(495), .W33TO42(256), .W33TO43(-991), .W33TO44(-825), .W33TO45(-957), .W33TO46(193), .W33TO47(93), .W33TO48(-497), .W33TO49(583), .W33TO50(-662), .W33TO51(-192), .W33TO52(-210), .W33TO53(737), .W33TO54(-999), .W33TO55(164), .W33TO56(349), .W33TO57(362), .W33TO58(-869), .W33TO59(-708), .W33TO60(155), .W33TO61(428), .W33TO62(-575), .W33TO63(660), .W34TO0(-625), .W34TO1(-534), .W34TO2(-840), .W34TO3(-632), .W34TO4(-167), .W34TO5(-671), .W34TO6(140), .W34TO7(486), .W34TO8(-368), .W34TO9(-10), .W34TO10(-197), .W34TO11(-743), .W34TO12(-818), .W34TO13(771), .W34TO14(-926), .W34TO15(23), .W34TO16(-460), .W34TO17(773), .W34TO18(-248), .W34TO19(-594), .W34TO20(652), .W34TO21(-139), .W34TO22(-533), .W34TO23(184), .W34TO24(-633), .W34TO25(787), .W34TO26(117), .W34TO27(-99), .W34TO28(-617), .W34TO29(-662), .W34TO30(-405), .W34TO31(-374), .W34TO32(26), .W34TO33(-540), .W34TO34(169), .W34TO35(735), .W34TO36(-708), .W34TO37(530), .W34TO38(208), .W34TO39(-293), .W34TO40(157), .W34TO41(645), .W34TO42(-891), .W34TO43(419), .W34TO44(790), .W34TO45(-499), .W34TO46(-385), .W34TO47(-881), .W34TO48(-745), .W34TO49(201), .W34TO50(855), .W34TO51(-678), .W34TO52(480), .W34TO53(84), .W34TO54(-468), .W34TO55(-140), .W34TO56(79), .W34TO57(375), .W34TO58(-488), .W34TO59(-48), .W34TO60(781), .W34TO61(-656), .W34TO62(-142), .W34TO63(487), .W35TO0(521), .W35TO1(-203), .W35TO2(-233), .W35TO3(-43), .W35TO4(-437), .W35TO5(178), .W35TO6(249), .W35TO7(-99), .W35TO8(-112), .W35TO9(-789), .W35TO10(698), .W35TO11(258), .W35TO12(-581), .W35TO13(910), .W35TO14(315), .W35TO15(180), .W35TO16(126), .W35TO17(796), .W35TO18(930), .W35TO19(-507), .W35TO20(350), .W35TO21(-816), .W35TO22(138), .W35TO23(528), .W35TO24(-544), .W35TO25(493), .W35TO26(997), .W35TO27(-376), .W35TO28(-80), .W35TO29(952), .W35TO30(688), .W35TO31(558), .W35TO32(327), .W35TO33(-594), .W35TO34(250), .W35TO35(0), .W35TO36(-487), .W35TO37(-395), .W35TO38(-191), .W35TO39(-847), .W35TO40(-932), .W35TO41(754), .W35TO42(371), .W35TO43(-494), .W35TO44(-484), .W35TO45(208), .W35TO46(-352), .W35TO47(91), .W35TO48(-517), .W35TO49(727), .W35TO50(778), .W35TO51(406), .W35TO52(-82), .W35TO53(458), .W35TO54(-545), .W35TO55(523), .W35TO56(500), .W35TO57(78), .W35TO58(885), .W35TO59(137), .W35TO60(-47), .W35TO61(495), .W35TO62(674), .W35TO63(-299), .W36TO0(68), .W36TO1(-434), .W36TO2(-573), .W36TO3(540), .W36TO4(-245), .W36TO5(-534), .W36TO6(969), .W36TO7(-119), .W36TO8(-883), .W36TO9(424), .W36TO10(-843), .W36TO11(134), .W36TO12(297), .W36TO13(149), .W36TO14(59), .W36TO15(4), .W36TO16(-584), .W36TO17(301), .W36TO18(-698), .W36TO19(-762), .W36TO20(-685), .W36TO21(395), .W36TO22(-578), .W36TO23(-35), .W36TO24(-853), .W36TO25(922), .W36TO26(-468), .W36TO27(647), .W36TO28(754), .W36TO29(-274), .W36TO30(665), .W36TO31(-219), .W36TO32(-622), .W36TO33(664), .W36TO34(-461), .W36TO35(261), .W36TO36(198), .W36TO37(726), .W36TO38(-816), .W36TO39(-344), .W36TO40(365), .W36TO41(-260), .W36TO42(136), .W36TO43(-854), .W36TO44(-88), .W36TO45(-829), .W36TO46(884), .W36TO47(628), .W36TO48(-818), .W36TO49(93), .W36TO50(-995), .W36TO51(572), .W36TO52(275), .W36TO53(678), .W36TO54(-608), .W36TO55(-203), .W36TO56(441), .W36TO57(390), .W36TO58(-16), .W36TO59(-428), .W36TO60(349), .W36TO61(978), .W36TO62(-860), .W36TO63(93), .W37TO0(11), .W37TO1(456), .W37TO2(866), .W37TO3(-479), .W37TO4(-388), .W37TO5(470), .W37TO6(882), .W37TO7(217), .W37TO8(706), .W37TO9(-533), .W37TO10(450), .W37TO11(251), .W37TO12(350), .W37TO13(-809), .W37TO14(809), .W37TO15(165), .W37TO16(-341), .W37TO17(308), .W37TO18(-304), .W37TO19(-696), .W37TO20(-481), .W37TO21(-16), .W37TO22(475), .W37TO23(-507), .W37TO24(45), .W37TO25(894), .W37TO26(-870), .W37TO27(-948), .W37TO28(-236), .W37TO29(-599), .W37TO30(286), .W37TO31(-542), .W37TO32(239), .W37TO33(739), .W37TO34(-778), .W37TO35(22), .W37TO36(-941), .W37TO37(415), .W37TO38(-673), .W37TO39(261), .W37TO40(-924), .W37TO41(902), .W37TO42(-134), .W37TO43(-769), .W37TO44(353), .W37TO45(775), .W37TO46(-463), .W37TO47(-153), .W37TO48(728), .W37TO49(495), .W37TO50(-191), .W37TO51(-326), .W37TO52(-839), .W37TO53(56), .W37TO54(-958), .W37TO55(-374), .W37TO56(43), .W37TO57(398), .W37TO58(-832), .W37TO59(241), .W37TO60(-684), .W37TO61(930), .W37TO62(-741), .W37TO63(9), .W38TO0(-936), .W38TO1(-23), .W38TO2(-113), .W38TO3(-671), .W38TO4(-344), .W38TO5(818), .W38TO6(545), .W38TO7(-230), .W38TO8(-758), .W38TO9(-372), .W38TO10(-587), .W38TO11(-94), .W38TO12(-963), .W38TO13(-936), .W38TO14(-245), .W38TO15(245), .W38TO16(161), .W38TO17(-458), .W38TO18(594), .W38TO19(-250), .W38TO20(-233), .W38TO21(542), .W38TO22(-238), .W38TO23(663), .W38TO24(968), .W38TO25(-29), .W38TO26(8), .W38TO27(639), .W38TO28(-402), .W38TO29(-552), .W38TO30(-158), .W38TO31(590), .W38TO32(104), .W38TO33(670), .W38TO34(499), .W38TO35(512), .W38TO36(-99), .W38TO37(-485), .W38TO38(659), .W38TO39(844), .W38TO40(-896), .W38TO41(143), .W38TO42(-808), .W38TO43(390), .W38TO44(-755), .W38TO45(876), .W38TO46(-37), .W38TO47(476), .W38TO48(681), .W38TO49(-557), .W38TO50(-78), .W38TO51(-307), .W38TO52(-344), .W38TO53(614), .W38TO54(-653), .W38TO55(603), .W38TO56(-121), .W38TO57(187), .W38TO58(659), .W38TO59(747), .W38TO60(-844), .W38TO61(-969), .W38TO62(-986), .W38TO63(345), .W39TO0(-901), .W39TO1(714), .W39TO2(-228), .W39TO3(-245), .W39TO4(768), .W39TO5(419), .W39TO6(55), .W39TO7(-869), .W39TO8(81), .W39TO9(503), .W39TO10(421), .W39TO11(-924), .W39TO12(768), .W39TO13(318), .W39TO14(436), .W39TO15(611), .W39TO16(-344), .W39TO17(295), .W39TO18(-202), .W39TO19(-64), .W39TO20(452), .W39TO21(859), .W39TO22(-289), .W39TO23(394), .W39TO24(954), .W39TO25(805), .W39TO26(939), .W39TO27(-802), .W39TO28(-658), .W39TO29(432), .W39TO30(-19), .W39TO31(430), .W39TO32(464), .W39TO33(769), .W39TO34(-473), .W39TO35(-913), .W39TO36(-923), .W39TO37(813), .W39TO38(139), .W39TO39(869), .W39TO40(755), .W39TO41(542), .W39TO42(438), .W39TO43(-946), .W39TO44(-993), .W39TO45(972), .W39TO46(-567), .W39TO47(-747), .W39TO48(-54), .W39TO49(-292), .W39TO50(-690), .W39TO51(857), .W39TO52(46), .W39TO53(-43), .W39TO54(-741), .W39TO55(-673), .W39TO56(-197), .W39TO57(406), .W39TO58(-648), .W39TO59(862), .W39TO60(756), .W39TO61(-385), .W39TO62(490), .W39TO63(838), .W40TO0(-102), .W40TO1(-111), .W40TO2(-628), .W40TO3(-688), .W40TO4(-331), .W40TO5(-26), .W40TO6(-769), .W40TO7(93), .W40TO8(-449), .W40TO9(684), .W40TO10(274), .W40TO11(-144), .W40TO12(38), .W40TO13(675), .W40TO14(-182), .W40TO15(-636), .W40TO16(600), .W40TO17(-685), .W40TO18(651), .W40TO19(-822), .W40TO20(-313), .W40TO21(136), .W40TO22(726), .W40TO23(305), .W40TO24(-743), .W40TO25(726), .W40TO26(-770), .W40TO27(-757), .W40TO28(989), .W40TO29(-656), .W40TO30(-271), .W40TO31(138), .W40TO32(513), .W40TO33(-666), .W40TO34(837), .W40TO35(-14), .W40TO36(-606), .W40TO37(-64), .W40TO38(-706), .W40TO39(-651), .W40TO40(450), .W40TO41(-813), .W40TO42(-681), .W40TO43(-658), .W40TO44(346), .W40TO45(750), .W40TO46(9), .W40TO47(-495), .W40TO48(227), .W40TO49(752), .W40TO50(-943), .W40TO51(-547), .W40TO52(271), .W40TO53(620), .W40TO54(129), .W40TO55(-619), .W40TO56(208), .W40TO57(535), .W40TO58(-491), .W40TO59(-10), .W40TO60(199), .W40TO61(562), .W40TO62(434), .W40TO63(-256), .W41TO0(-688), .W41TO1(-142), .W41TO2(-563), .W41TO3(-668), .W41TO4(-648), .W41TO5(-516), .W41TO6(755), .W41TO7(116), .W41TO8(-315), .W41TO9(-334), .W41TO10(160), .W41TO11(-784), .W41TO12(606), .W41TO13(628), .W41TO14(800), .W41TO15(416), .W41TO16(106), .W41TO17(908), .W41TO18(260), .W41TO19(-865), .W41TO20(817), .W41TO21(505), .W41TO22(-595), .W41TO23(78), .W41TO24(952), .W41TO25(187), .W41TO26(873), .W41TO27(-506), .W41TO28(405), .W41TO29(-846), .W41TO30(583), .W41TO31(-965), .W41TO32(-134), .W41TO33(763), .W41TO34(-191), .W41TO35(891), .W41TO36(183), .W41TO37(-231), .W41TO38(503), .W41TO39(-796), .W41TO40(-467), .W41TO41(-890), .W41TO42(109), .W41TO43(122), .W41TO44(814), .W41TO45(85), .W41TO46(389), .W41TO47(-377), .W41TO48(-58), .W41TO49(-308), .W41TO50(-595), .W41TO51(-544), .W41TO52(-571), .W41TO53(865), .W41TO54(994), .W41TO55(-40), .W41TO56(581), .W41TO57(-119), .W41TO58(-496), .W41TO59(-896), .W41TO60(954), .W41TO61(366), .W41TO62(-28), .W41TO63(691), .W42TO0(415), .W42TO1(274), .W42TO2(-295), .W42TO3(-170), .W42TO4(403), .W42TO5(33), .W42TO6(-844), .W42TO7(576), .W42TO8(651), .W42TO9(546), .W42TO10(650), .W42TO11(-253), .W42TO12(198), .W42TO13(-468), .W42TO14(-644), .W42TO15(-514), .W42TO16(754), .W42TO17(-616), .W42TO18(507), .W42TO19(126), .W42TO20(876), .W42TO21(927), .W42TO22(911), .W42TO23(-598), .W42TO24(787), .W42TO25(-857), .W42TO26(-327), .W42TO27(-907), .W42TO28(-68), .W42TO29(447), .W42TO30(984), .W42TO31(-394), .W42TO32(-709), .W42TO33(616), .W42TO34(-798), .W42TO35(173), .W42TO36(-870), .W42TO37(-273), .W42TO38(407), .W42TO39(-774), .W42TO40(192), .W42TO41(-611), .W42TO42(535), .W42TO43(784), .W42TO44(393), .W42TO45(518), .W42TO46(-199), .W42TO47(-353), .W42TO48(41), .W42TO49(295), .W42TO50(-610), .W42TO51(-353), .W42TO52(354), .W42TO53(-900), .W42TO54(-883), .W42TO55(351), .W42TO56(690), .W42TO57(342), .W42TO58(18), .W42TO59(-524), .W42TO60(-672), .W42TO61(-690), .W42TO62(-493), .W42TO63(71), .W43TO0(963), .W43TO1(-693), .W43TO2(187), .W43TO3(475), .W43TO4(808), .W43TO5(-799), .W43TO6(-26), .W43TO7(246), .W43TO8(845), .W43TO9(-424), .W43TO10(-138), .W43TO11(-989), .W43TO12(217), .W43TO13(396), .W43TO14(-494), .W43TO15(918), .W43TO16(187), .W43TO17(-927), .W43TO18(-28), .W43TO19(283), .W43TO20(-176), .W43TO21(-58), .W43TO22(899), .W43TO23(-651), .W43TO24(468), .W43TO25(-39), .W43TO26(436), .W43TO27(-32), .W43TO28(-448), .W43TO29(-601), .W43TO30(791), .W43TO31(832), .W43TO32(431), .W43TO33(199), .W43TO34(-618), .W43TO35(75), .W43TO36(-850), .W43TO37(-343), .W43TO38(533), .W43TO39(356), .W43TO40(-800), .W43TO41(-618), .W43TO42(-583), .W43TO43(725), .W43TO44(788), .W43TO45(-570), .W43TO46(-257), .W43TO47(239), .W43TO48(-345), .W43TO49(747), .W43TO50(-660), .W43TO51(369), .W43TO52(-727), .W43TO53(-531), .W43TO54(46), .W43TO55(772), .W43TO56(638), .W43TO57(-429), .W43TO58(356), .W43TO59(-773), .W43TO60(-68), .W43TO61(566), .W43TO62(771), .W43TO63(949), .W44TO0(692), .W44TO1(243), .W44TO2(677), .W44TO3(-502), .W44TO4(223), .W44TO5(-104), .W44TO6(-681), .W44TO7(-222), .W44TO8(-734), .W44TO9(824), .W44TO10(-377), .W44TO11(-942), .W44TO12(-339), .W44TO13(-525), .W44TO14(-422), .W44TO15(-872), .W44TO16(-837), .W44TO17(290), .W44TO18(213), .W44TO19(270), .W44TO20(-307), .W44TO21(31), .W44TO22(471), .W44TO23(241), .W44TO24(358), .W44TO25(944), .W44TO26(-467), .W44TO27(-819), .W44TO28(132), .W44TO29(700), .W44TO30(942), .W44TO31(-153), .W44TO32(-658), .W44TO33(-641), .W44TO34(-934), .W44TO35(-799), .W44TO36(592), .W44TO37(-580), .W44TO38(-215), .W44TO39(-952), .W44TO40(-874), .W44TO41(191), .W44TO42(-250), .W44TO43(-238), .W44TO44(599), .W44TO45(-363), .W44TO46(261), .W44TO47(679), .W44TO48(-33), .W44TO49(-291), .W44TO50(-125), .W44TO51(774), .W44TO52(741), .W44TO53(-356), .W44TO54(452), .W44TO55(-36), .W44TO56(63), .W44TO57(461), .W44TO58(485), .W44TO59(-105), .W44TO60(195), .W44TO61(-507), .W44TO62(195), .W44TO63(-222), .W45TO0(-905), .W45TO1(563), .W45TO2(-876), .W45TO3(117), .W45TO4(-216), .W45TO5(-915), .W45TO6(-884), .W45TO7(-836), .W45TO8(625), .W45TO9(-5), .W45TO10(7), .W45TO11(-937), .W45TO12(965), .W45TO13(-846), .W45TO14(960), .W45TO15(138), .W45TO16(-894), .W45TO17(924), .W45TO18(826), .W45TO19(976), .W45TO20(832), .W45TO21(963), .W45TO22(-751), .W45TO23(-626), .W45TO24(169), .W45TO25(-862), .W45TO26(639), .W45TO27(-547), .W45TO28(-241), .W45TO29(-114), .W45TO30(520), .W45TO31(309), .W45TO32(42), .W45TO33(892), .W45TO34(108), .W45TO35(530), .W45TO36(-113), .W45TO37(-299), .W45TO38(-793), .W45TO39(-789), .W45TO40(81), .W45TO41(-504), .W45TO42(-968), .W45TO43(-632), .W45TO44(277), .W45TO45(-806), .W45TO46(601), .W45TO47(-979), .W45TO48(-498), .W45TO49(445), .W45TO50(-789), .W45TO51(804), .W45TO52(444), .W45TO53(769), .W45TO54(-618), .W45TO55(-28), .W45TO56(779), .W45TO57(-446), .W45TO58(-517), .W45TO59(58), .W45TO60(778), .W45TO61(982), .W45TO62(-203), .W45TO63(-401), .W46TO0(156), .W46TO1(794), .W46TO2(-603), .W46TO3(823), .W46TO4(-778), .W46TO5(688), .W46TO6(-816), .W46TO7(-636), .W46TO8(839), .W46TO9(566), .W46TO10(-958), .W46TO11(477), .W46TO12(-910), .W46TO13(-96), .W46TO14(414), .W46TO15(-97), .W46TO16(957), .W46TO17(-753), .W46TO18(-549), .W46TO19(-749), .W46TO20(-609), .W46TO21(-764), .W46TO22(-353), .W46TO23(964), .W46TO24(-887), .W46TO25(50), .W46TO26(653), .W46TO27(923), .W46TO28(268), .W46TO29(632), .W46TO30(950), .W46TO31(626), .W46TO32(234), .W46TO33(3), .W46TO34(-573), .W46TO35(-672), .W46TO36(-70), .W46TO37(733), .W46TO38(-941), .W46TO39(871), .W46TO40(740), .W46TO41(-535), .W46TO42(679), .W46TO43(-22), .W46TO44(543), .W46TO45(358), .W46TO46(-194), .W46TO47(144), .W46TO48(71), .W46TO49(724), .W46TO50(256), .W46TO51(126), .W46TO52(885), .W46TO53(-978), .W46TO54(526), .W46TO55(564), .W46TO56(-805), .W46TO57(470), .W46TO58(699), .W46TO59(713), .W46TO60(-441), .W46TO61(450), .W46TO62(-524), .W46TO63(-972), .W47TO0(849), .W47TO1(-132), .W47TO2(382), .W47TO3(190), .W47TO4(-360), .W47TO5(969), .W47TO6(-934), .W47TO7(473), .W47TO8(-887), .W47TO9(-572), .W47TO10(-169), .W47TO11(-70), .W47TO12(631), .W47TO13(-918), .W47TO14(-979), .W47TO15(-445), .W47TO16(125), .W47TO17(947), .W47TO18(866), .W47TO19(-59), .W47TO20(-910), .W47TO21(-134), .W47TO22(595), .W47TO23(699), .W47TO24(-321), .W47TO25(411), .W47TO26(971), .W47TO27(871), .W47TO28(-299), .W47TO29(765), .W47TO30(433), .W47TO31(741), .W47TO32(-35), .W47TO33(984), .W47TO34(-553), .W47TO35(-506), .W47TO36(854), .W47TO37(864), .W47TO38(-540), .W47TO39(697), .W47TO40(210), .W47TO41(-624), .W47TO42(99), .W47TO43(641), .W47TO44(-253), .W47TO45(220), .W47TO46(-461), .W47TO47(-753), .W47TO48(503), .W47TO49(-953), .W47TO50(-214), .W47TO51(-467), .W47TO52(818), .W47TO53(-394), .W47TO54(71), .W47TO55(-483), .W47TO56(341), .W47TO57(803), .W47TO58(92), .W47TO59(442), .W47TO60(465), .W47TO61(-418), .W47TO62(-393), .W47TO63(775), .W48TO0(-892), .W48TO1(-471), .W48TO2(-78), .W48TO3(-566), .W48TO4(275), .W48TO5(843), .W48TO6(765), .W48TO7(254), .W48TO8(844), .W48TO9(163), .W48TO10(490), .W48TO11(287), .W48TO12(21), .W48TO13(451), .W48TO14(-613), .W48TO15(724), .W48TO16(-637), .W48TO17(-354), .W48TO18(-125), .W48TO19(-342), .W48TO20(-81), .W48TO21(-326), .W48TO22(766), .W48TO23(-428), .W48TO24(249), .W48TO25(-701), .W48TO26(-362), .W48TO27(820), .W48TO28(-195), .W48TO29(-611), .W48TO30(-839), .W48TO31(14), .W48TO32(-40), .W48TO33(584), .W48TO34(-437), .W48TO35(301), .W48TO36(40), .W48TO37(-537), .W48TO38(-727), .W48TO39(-609), .W48TO40(602), .W48TO41(246), .W48TO42(-942), .W48TO43(593), .W48TO44(-474), .W48TO45(433), .W48TO46(664), .W48TO47(-962), .W48TO48(-73), .W48TO49(-385), .W48TO50(669), .W48TO51(-737), .W48TO52(855), .W48TO53(-939), .W48TO54(679), .W48TO55(558), .W48TO56(-143), .W48TO57(-745), .W48TO58(-196), .W48TO59(472), .W48TO60(-491), .W48TO61(973), .W48TO62(-339), .W48TO63(-906), .W49TO0(52), .W49TO1(8), .W49TO2(-145), .W49TO3(-388), .W49TO4(944), .W49TO5(331), .W49TO6(44), .W49TO7(660), .W49TO8(366), .W49TO9(-317), .W49TO10(-209), .W49TO11(231), .W49TO12(875), .W49TO13(-25), .W49TO14(-156), .W49TO15(-302), .W49TO16(-770), .W49TO17(-785), .W49TO18(-989), .W49TO19(532), .W49TO20(-323), .W49TO21(-213), .W49TO22(-685), .W49TO23(710), .W49TO24(832), .W49TO25(-779), .W49TO26(-879), .W49TO27(344), .W49TO28(688), .W49TO29(809), .W49TO30(240), .W49TO31(-733), .W49TO32(715), .W49TO33(-636), .W49TO34(-406), .W49TO35(720), .W49TO36(528), .W49TO37(820), .W49TO38(-861), .W49TO39(278), .W49TO40(-381), .W49TO41(993), .W49TO42(-247), .W49TO43(-681), .W49TO44(-102), .W49TO45(-24), .W49TO46(-705), .W49TO47(-456), .W49TO48(157), .W49TO49(951), .W49TO50(816), .W49TO51(454), .W49TO52(-625), .W49TO53(352), .W49TO54(-648), .W49TO55(15), .W49TO56(-671), .W49TO57(664), .W49TO58(971), .W49TO59(-993), .W49TO60(-114), .W49TO61(-852), .W49TO62(-146), .W49TO63(-830), .W50TO0(-522), .W50TO1(720), .W50TO2(442), .W50TO3(-271), .W50TO4(-781), .W50TO5(75), .W50TO6(608), .W50TO7(346), .W50TO8(-25), .W50TO9(-678), .W50TO10(-963), .W50TO11(-556), .W50TO12(708), .W50TO13(-496), .W50TO14(-517), .W50TO15(506), .W50TO16(157), .W50TO17(-746), .W50TO18(380), .W50TO19(949), .W50TO20(801), .W50TO21(-758), .W50TO22(342), .W50TO23(-63), .W50TO24(121), .W50TO25(116), .W50TO26(-818), .W50TO27(-507), .W50TO28(558), .W50TO29(28), .W50TO30(174), .W50TO31(974), .W50TO32(377), .W50TO33(-956), .W50TO34(417), .W50TO35(-67), .W50TO36(-59), .W50TO37(-489), .W50TO38(545), .W50TO39(-408), .W50TO40(-320), .W50TO41(-81), .W50TO42(-22), .W50TO43(430), .W50TO44(-793), .W50TO45(-477), .W50TO46(332), .W50TO47(298), .W50TO48(-21), .W50TO49(459), .W50TO50(60), .W50TO51(181), .W50TO52(-390), .W50TO53(106), .W50TO54(11), .W50TO55(-997), .W50TO56(-556), .W50TO57(-294), .W50TO58(-155), .W50TO59(-641), .W50TO60(-487), .W50TO61(713), .W50TO62(615), .W50TO63(450), .W51TO0(-848), .W51TO1(759), .W51TO2(706), .W51TO3(-597), .W51TO4(-501), .W51TO5(860), .W51TO6(403), .W51TO7(64), .W51TO8(-493), .W51TO9(134), .W51TO10(-189), .W51TO11(-371), .W51TO12(-384), .W51TO13(-306), .W51TO14(74), .W51TO15(-761), .W51TO16(467), .W51TO17(630), .W51TO18(63), .W51TO19(-781), .W51TO20(480), .W51TO21(531), .W51TO22(715), .W51TO23(215), .W51TO24(564), .W51TO25(-180), .W51TO26(889), .W51TO27(-524), .W51TO28(-408), .W51TO29(-629), .W51TO30(786), .W51TO31(-484), .W51TO32(132), .W51TO33(479), .W51TO34(870), .W51TO35(309), .W51TO36(318), .W51TO37(-943), .W51TO38(359), .W51TO39(271), .W51TO40(-695), .W51TO41(531), .W51TO42(-438), .W51TO43(-46), .W51TO44(-463), .W51TO45(771), .W51TO46(918), .W51TO47(-510), .W51TO48(921), .W51TO49(-39), .W51TO50(352), .W51TO51(715), .W51TO52(-731), .W51TO53(-217), .W51TO54(-255), .W51TO55(899), .W51TO56(-474), .W51TO57(814), .W51TO58(-904), .W51TO59(-928), .W51TO60(535), .W51TO61(-210), .W51TO62(-57), .W51TO63(248), .W52TO0(727), .W52TO1(920), .W52TO2(-754), .W52TO3(-767), .W52TO4(-887), .W52TO5(-586), .W52TO6(956), .W52TO7(-606), .W52TO8(244), .W52TO9(-497), .W52TO10(-52), .W52TO11(-395), .W52TO12(294), .W52TO13(845), .W52TO14(-232), .W52TO15(570), .W52TO16(238), .W52TO17(-323), .W52TO18(763), .W52TO19(-845), .W52TO20(45), .W52TO21(-545), .W52TO22(-446), .W52TO23(343), .W52TO24(700), .W52TO25(749), .W52TO26(787), .W52TO27(952), .W52TO28(458), .W52TO29(-598), .W52TO30(-748), .W52TO31(56), .W52TO32(234), .W52TO33(66), .W52TO34(911), .W52TO35(746), .W52TO36(-558), .W52TO37(36), .W52TO38(389), .W52TO39(472), .W52TO40(85), .W52TO41(-278), .W52TO42(820), .W52TO43(420), .W52TO44(988), .W52TO45(-278), .W52TO46(504), .W52TO47(-769), .W52TO48(-968), .W52TO49(-611), .W52TO50(-683), .W52TO51(-275), .W52TO52(346), .W52TO53(82), .W52TO54(-594), .W52TO55(-33), .W52TO56(521), .W52TO57(783), .W52TO58(746), .W52TO59(-527), .W52TO60(-160), .W52TO61(485), .W52TO62(778), .W52TO63(176), .W53TO0(307), .W53TO1(387), .W53TO2(-664), .W53TO3(-333), .W53TO4(-407), .W53TO5(-989), .W53TO6(987), .W53TO7(219), .W53TO8(917), .W53TO9(924), .W53TO10(-745), .W53TO11(263), .W53TO12(162), .W53TO13(-72), .W53TO14(131), .W53TO15(72), .W53TO16(-392), .W53TO17(906), .W53TO18(-949), .W53TO19(822), .W53TO20(111), .W53TO21(610), .W53TO22(-830), .W53TO23(-862), .W53TO24(-976), .W53TO25(265), .W53TO26(564), .W53TO27(799), .W53TO28(-155), .W53TO29(339), .W53TO30(16), .W53TO31(235), .W53TO32(-147), .W53TO33(-457), .W53TO34(900), .W53TO35(-178), .W53TO36(-344), .W53TO37(-194), .W53TO38(521), .W53TO39(977), .W53TO40(652), .W53TO41(914), .W53TO42(2), .W53TO43(-981), .W53TO44(-41), .W53TO45(-946), .W53TO46(879), .W53TO47(-48), .W53TO48(904), .W53TO49(313), .W53TO50(962), .W53TO51(-716), .W53TO52(567), .W53TO53(714), .W53TO54(-604), .W53TO55(524), .W53TO56(-757), .W53TO57(98), .W53TO58(-188), .W53TO59(-402), .W53TO60(704), .W53TO61(759), .W53TO62(318), .W53TO63(-178), .W54TO0(-718), .W54TO1(-407), .W54TO2(854), .W54TO3(-93), .W54TO4(-52), .W54TO5(619), .W54TO6(-563), .W54TO7(290), .W54TO8(876), .W54TO9(-43), .W54TO10(572), .W54TO11(-314), .W54TO12(-6), .W54TO13(781), .W54TO14(-565), .W54TO15(981), .W54TO16(-821), .W54TO17(577), .W54TO18(681), .W54TO19(355), .W54TO20(925), .W54TO21(-40), .W54TO22(436), .W54TO23(362), .W54TO24(-688), .W54TO25(805), .W54TO26(516), .W54TO27(859), .W54TO28(243), .W54TO29(-946), .W54TO30(265), .W54TO31(-318), .W54TO32(191), .W54TO33(283), .W54TO34(-308), .W54TO35(418), .W54TO36(-669), .W54TO37(400), .W54TO38(222), .W54TO39(-663), .W54TO40(758), .W54TO41(-265), .W54TO42(922), .W54TO43(-333), .W54TO44(-431), .W54TO45(-399), .W54TO46(806), .W54TO47(-558), .W54TO48(-975), .W54TO49(334), .W54TO50(539), .W54TO51(190), .W54TO52(626), .W54TO53(150), .W54TO54(-237), .W54TO55(-766), .W54TO56(16), .W54TO57(537), .W54TO58(-949), .W54TO59(570), .W54TO60(265), .W54TO61(-592), .W54TO62(-632), .W54TO63(432), .W55TO0(624), .W55TO1(-857), .W55TO2(986), .W55TO3(506), .W55TO4(129), .W55TO5(-409), .W55TO6(-288), .W55TO7(-176), .W55TO8(-269), .W55TO9(-15), .W55TO10(353), .W55TO11(839), .W55TO12(586), .W55TO13(-71), .W55TO14(413), .W55TO15(879), .W55TO16(842), .W55TO17(189), .W55TO18(905), .W55TO19(395), .W55TO20(591), .W55TO21(149), .W55TO22(132), .W55TO23(584), .W55TO24(972), .W55TO25(-916), .W55TO26(-107), .W55TO27(-927), .W55TO28(821), .W55TO29(133), .W55TO30(-844), .W55TO31(-390), .W55TO32(-389), .W55TO33(966), .W55TO34(-253), .W55TO35(209), .W55TO36(-803), .W55TO37(-123), .W55TO38(-285), .W55TO39(-324), .W55TO40(-857), .W55TO41(973), .W55TO42(-427), .W55TO43(521), .W55TO44(-29), .W55TO45(-968), .W55TO46(-764), .W55TO47(-542), .W55TO48(-461), .W55TO49(699), .W55TO50(-502), .W55TO51(300), .W55TO52(592), .W55TO53(-469), .W55TO54(-269), .W55TO55(90), .W55TO56(802), .W55TO57(374), .W55TO58(-888), .W55TO59(975), .W55TO60(-930), .W55TO61(655), .W55TO62(-771), .W55TO63(723), .W56TO0(-457), .W56TO1(-418), .W56TO2(-590), .W56TO3(905), .W56TO4(-966), .W56TO5(557), .W56TO6(274), .W56TO7(740), .W56TO8(36), .W56TO9(-40), .W56TO10(-972), .W56TO11(295), .W56TO12(161), .W56TO13(223), .W56TO14(-396), .W56TO15(717), .W56TO16(13), .W56TO17(136), .W56TO18(711), .W56TO19(-364), .W56TO20(115), .W56TO21(-463), .W56TO22(-286), .W56TO23(596), .W56TO24(364), .W56TO25(-914), .W56TO26(-14), .W56TO27(-876), .W56TO28(-591), .W56TO29(201), .W56TO30(-114), .W56TO31(-486), .W56TO32(41), .W56TO33(-234), .W56TO34(-497), .W56TO35(192), .W56TO36(771), .W56TO37(-505), .W56TO38(-424), .W56TO39(-602), .W56TO40(-599), .W56TO41(-195), .W56TO42(893), .W56TO43(-605), .W56TO44(-884), .W56TO45(-82), .W56TO46(793), .W56TO47(-812), .W56TO48(173), .W56TO49(962), .W56TO50(-607), .W56TO51(407), .W56TO52(-438), .W56TO53(746), .W56TO54(352), .W56TO55(398), .W56TO56(302), .W56TO57(-985), .W56TO58(791), .W56TO59(925), .W56TO60(550), .W56TO61(344), .W56TO62(45), .W56TO63(483), .W57TO0(-804), .W57TO1(-967), .W57TO2(961), .W57TO3(-67), .W57TO4(-606), .W57TO5(522), .W57TO6(-981), .W57TO7(-876), .W57TO8(99), .W57TO9(874), .W57TO10(739), .W57TO11(812), .W57TO12(-624), .W57TO13(920), .W57TO14(-813), .W57TO15(-735), .W57TO16(354), .W57TO17(904), .W57TO18(49), .W57TO19(-103), .W57TO20(-485), .W57TO21(963), .W57TO22(129), .W57TO23(-839), .W57TO24(-128), .W57TO25(58), .W57TO26(-994), .W57TO27(-84), .W57TO28(411), .W57TO29(32), .W57TO30(-430), .W57TO31(399), .W57TO32(808), .W57TO33(947), .W57TO34(-873), .W57TO35(98), .W57TO36(89), .W57TO37(681), .W57TO38(662), .W57TO39(-9), .W57TO40(-438), .W57TO41(585), .W57TO42(345), .W57TO43(-250), .W57TO44(-889), .W57TO45(892), .W57TO46(-299), .W57TO47(62), .W57TO48(-146), .W57TO49(60), .W57TO50(-836), .W57TO51(-319), .W57TO52(-947), .W57TO53(-661), .W57TO54(287), .W57TO55(883), .W57TO56(344), .W57TO57(-38), .W57TO58(790), .W57TO59(-26), .W57TO60(-742), .W57TO61(-574), .W57TO62(178), .W57TO63(-112), .W58TO0(-621), .W58TO1(392), .W58TO2(-286), .W58TO3(-12), .W58TO4(657), .W58TO5(272), .W58TO6(729), .W58TO7(-314), .W58TO8(840), .W58TO9(-622), .W58TO10(-393), .W58TO11(-690), .W58TO12(-584), .W58TO13(-305), .W58TO14(-529), .W58TO15(-162), .W58TO16(620), .W58TO17(-927), .W58TO18(-201), .W58TO19(-989), .W58TO20(793), .W58TO21(272), .W58TO22(149), .W58TO23(639), .W58TO24(945), .W58TO25(849), .W58TO26(-42), .W58TO27(635), .W58TO28(-59), .W58TO29(-65), .W58TO30(437), .W58TO31(510), .W58TO32(720), .W58TO33(-62), .W58TO34(297), .W58TO35(132), .W58TO36(475), .W58TO37(69), .W58TO38(198), .W58TO39(-727), .W58TO40(-67), .W58TO41(-208), .W58TO42(-722), .W58TO43(-206), .W58TO44(227), .W58TO45(-732), .W58TO46(741), .W58TO47(90), .W58TO48(311), .W58TO49(-87), .W58TO50(308), .W58TO51(-747), .W58TO52(-545), .W58TO53(-757), .W58TO54(373), .W58TO55(-502), .W58TO56(-88), .W58TO57(-178), .W58TO58(994), .W58TO59(750), .W58TO60(-419), .W58TO61(805), .W58TO62(287), .W58TO63(261), .W59TO0(-322), .W59TO1(783), .W59TO2(505), .W59TO3(-760), .W59TO4(268), .W59TO5(-834), .W59TO6(652), .W59TO7(889), .W59TO8(-791), .W59TO9(-710), .W59TO10(-433), .W59TO11(-223), .W59TO12(-544), .W59TO13(645), .W59TO14(-172), .W59TO15(932), .W59TO16(-860), .W59TO17(974), .W59TO18(259), .W59TO19(-297), .W59TO20(-660), .W59TO21(-88), .W59TO22(-83), .W59TO23(409), .W59TO24(836), .W59TO25(-747), .W59TO26(-92), .W59TO27(329), .W59TO28(140), .W59TO29(202), .W59TO30(-775), .W59TO31(970), .W59TO32(-24), .W59TO33(-785), .W59TO34(-768), .W59TO35(206), .W59TO36(-888), .W59TO37(220), .W59TO38(-811), .W59TO39(754), .W59TO40(459), .W59TO41(558), .W59TO42(-296), .W59TO43(404), .W59TO44(113), .W59TO45(-73), .W59TO46(370), .W59TO47(-878), .W59TO48(-115), .W59TO49(-516), .W59TO50(-824), .W59TO51(-495), .W59TO52(-998), .W59TO53(986), .W59TO54(104), .W59TO55(511), .W59TO56(-872), .W59TO57(-707), .W59TO58(467), .W59TO59(649), .W59TO60(641), .W59TO61(-80), .W59TO62(-768), .W59TO63(399), .W60TO0(-84), .W60TO1(-217), .W60TO2(-732), .W60TO3(-818), .W60TO4(449), .W60TO5(576), .W60TO6(606), .W60TO7(888), .W60TO8(-476), .W60TO9(-817), .W60TO10(519), .W60TO11(-304), .W60TO12(-984), .W60TO13(-418), .W60TO14(280), .W60TO15(-567), .W60TO16(-195), .W60TO17(-977), .W60TO18(-952), .W60TO19(491), .W60TO20(192), .W60TO21(344), .W60TO22(-468), .W60TO23(-528), .W60TO24(528), .W60TO25(-344), .W60TO26(763), .W60TO27(-728), .W60TO28(-970), .W60TO29(-34), .W60TO30(780), .W60TO31(386), .W60TO32(-669), .W60TO33(-750), .W60TO34(511), .W60TO35(125), .W60TO36(72), .W60TO37(-926), .W60TO38(168), .W60TO39(-450), .W60TO40(710), .W60TO41(-638), .W60TO42(-777), .W60TO43(-665), .W60TO44(722), .W60TO45(436), .W60TO46(150), .W60TO47(-221), .W60TO48(-766), .W60TO49(140), .W60TO50(-260), .W60TO51(-792), .W60TO52(-494), .W60TO53(-799), .W60TO54(-830), .W60TO55(-310), .W60TO56(955), .W60TO57(112), .W60TO58(485), .W60TO59(652), .W60TO60(-204), .W60TO61(651), .W60TO62(11), .W60TO63(824), .W61TO0(529), .W61TO1(652), .W61TO2(361), .W61TO3(669), .W61TO4(720), .W61TO5(170), .W61TO6(619), .W61TO7(741), .W61TO8(546), .W61TO9(821), .W61TO10(-585), .W61TO11(219), .W61TO12(-994), .W61TO13(73), .W61TO14(635), .W61TO15(593), .W61TO16(-160), .W61TO17(-234), .W61TO18(707), .W61TO19(-157), .W61TO20(331), .W61TO21(602), .W61TO22(-539), .W61TO23(248), .W61TO24(-565), .W61TO25(-92), .W61TO26(48), .W61TO27(904), .W61TO28(938), .W61TO29(-493), .W61TO30(409), .W61TO31(622), .W61TO32(-623), .W61TO33(513), .W61TO34(-77), .W61TO35(-19), .W61TO36(306), .W61TO37(466), .W61TO38(-505), .W61TO39(-497), .W61TO40(926), .W61TO41(865), .W61TO42(438), .W61TO43(-106), .W61TO44(-203), .W61TO45(68), .W61TO46(-990), .W61TO47(372), .W61TO48(322), .W61TO49(814), .W61TO50(-726), .W61TO51(-656), .W61TO52(-709), .W61TO53(651), .W61TO54(39), .W61TO55(979), .W61TO56(-578), .W61TO57(237), .W61TO58(465), .W61TO59(-233), .W61TO60(-876), .W61TO61(-192), .W61TO62(-558), .W61TO63(-34), .W62TO0(-326), .W62TO1(493), .W62TO2(643), .W62TO3(706), .W62TO4(486), .W62TO5(123), .W62TO6(664), .W62TO7(431), .W62TO8(234), .W62TO9(938), .W62TO10(-918), .W62TO11(-450), .W62TO12(589), .W62TO13(-765), .W62TO14(-640), .W62TO15(672), .W62TO16(-320), .W62TO17(-384), .W62TO18(-102), .W62TO19(-211), .W62TO20(932), .W62TO21(-660), .W62TO22(-700), .W62TO23(-962), .W62TO24(624), .W62TO25(-711), .W62TO26(-947), .W62TO27(322), .W62TO28(-760), .W62TO29(-723), .W62TO30(-103), .W62TO31(-154), .W62TO32(242), .W62TO33(-452), .W62TO34(935), .W62TO35(-539), .W62TO36(-211), .W62TO37(-816), .W62TO38(-664), .W62TO39(-936), .W62TO40(313), .W62TO41(-91), .W62TO42(600), .W62TO43(-217), .W62TO44(-985), .W62TO45(607), .W62TO46(-946), .W62TO47(-365), .W62TO48(597), .W62TO49(197), .W62TO50(720), .W62TO51(478), .W62TO52(-897), .W62TO53(273), .W62TO54(-369), .W62TO55(822), .W62TO56(-88), .W62TO57(768), .W62TO58(-493), .W62TO59(55), .W62TO60(-912), .W62TO61(-594), .W62TO62(947), .W62TO63(-948), .W63TO0(846), .W63TO1(700), .W63TO2(-501), .W63TO3(-998), .W63TO4(474), .W63TO5(732), .W63TO6(-618), .W63TO7(951), .W63TO8(877), .W63TO9(541), .W63TO10(-447), .W63TO11(726), .W63TO12(325), .W63TO13(768), .W63TO14(19), .W63TO15(709), .W63TO16(286), .W63TO17(-783), .W63TO18(-535), .W63TO19(7), .W63TO20(-400), .W63TO21(129), .W63TO22(-723), .W63TO23(-289), .W63TO24(502), .W63TO25(475), .W63TO26(251), .W63TO27(-469), .W63TO28(-880), .W63TO29(-124), .W63TO30(732), .W63TO31(646), .W63TO32(722), .W63TO33(-407), .W63TO34(869), .W63TO35(-189), .W63TO36(-976), .W63TO37(-325), .W63TO38(423), .W63TO39(-721), .W63TO40(803), .W63TO41(534), .W63TO42(664), .W63TO43(541), .W63TO44(-41), .W63TO45(634), .W63TO46(-950), .W63TO47(-160), .W63TO48(284), .W63TO49(963), .W63TO50(-972), .W63TO51(-335), .W63TO52(121), .W63TO53(93), .W63TO54(-95), .W63TO55(-252), .W63TO56(961), .W63TO57(796), .W63TO58(-492), .W63TO59(-835), .W63TO60(610), .W63TO61(625), .W63TO62(-591), .W63TO63(313), .W64TO0(-251), .W64TO1(-842), .W64TO2(796), .W64TO3(-962), .W64TO4(302), .W64TO5(492), .W64TO6(-622), .W64TO7(796), .W64TO8(558), .W64TO9(549), .W64TO10(-530), .W64TO11(-729), .W64TO12(992), .W64TO13(612), .W64TO14(-254), .W64TO15(-751), .W64TO16(708), .W64TO17(-834), .W64TO18(-666), .W64TO19(-754), .W64TO20(-600), .W64TO21(-72), .W64TO22(-663), .W64TO23(811), .W64TO24(-172), .W64TO25(-198), .W64TO26(-509), .W64TO27(33), .W64TO28(29), .W64TO29(932), .W64TO30(678), .W64TO31(544), .W64TO32(-346), .W64TO33(570), .W64TO34(162), .W64TO35(-57), .W64TO36(-429), .W64TO37(622), .W64TO38(434), .W64TO39(238), .W64TO40(-916), .W64TO41(291), .W64TO42(302), .W64TO43(-723), .W64TO44(-503), .W64TO45(784), .W64TO46(990), .W64TO47(56), .W64TO48(-780), .W64TO49(-102), .W64TO50(728), .W64TO51(215), .W64TO52(24), .W64TO53(890), .W64TO54(-526), .W64TO55(-938), .W64TO56(-829), .W64TO57(-932), .W64TO58(-985), .W64TO59(-671), .W64TO60(172), .W64TO61(232), .W64TO62(-186), .W64TO63(-692)) layer0(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out0(con0[0]), .out1(con0[1]), .out2(con0[2]), .out3(con0[3]), .out4(con0[4]), .out5(con0[5]), .out6(con0[6]), .out7(con0[7]), .out8(con0[8]), .out9(con0[9]), .out10(con0[10]), .out11(con0[11]), .out12(con0[12]), .out13(con0[13]), .out14(con0[14]), .out15(con0[15]), .out16(con0[16]), .out17(con0[17]), .out18(con0[18]), .out19(con0[19]), .out20(con0[20]), .out21(con0[21]), .out22(con0[22]), .out23(con0[23]), .out24(con0[24]), .out25(con0[25]), .out26(con0[26]), .out27(con0[27]), .out28(con0[28]), .out29(con0[29]), .out30(con0[30]), .out31(con0[31]), .out32(con0[32]), .out33(con0[33]), .out34(con0[34]), .out35(con0[35]), .out36(con0[36]), .out37(con0[37]), .out38(con0[38]), .out39(con0[39]), .out40(con0[40]), .out41(con0[41]), .out42(con0[42]), .out43(con0[43]), .out44(con0[44]), .out45(con0[45]), .out46(con0[46]), .out47(con0[47]), .out48(con0[48]), .out49(con0[49]), .out50(con0[50]), .out51(con0[51]), .out52(con0[52]), .out53(con0[53]), .out54(con0[54]), .out55(con0[55]), .out56(con0[56]), .out57(con0[57]), .out58(con0[58]), .out59(con0[59]), .out60(con0[60]), .out61(con0[61]), .out62(con0[62]), .out63(con0[63]));
layer64in1out #(.BIAS0(-917), .W0TO0(971), .W1TO0(-582), .W2TO0(-107), .W3TO0(-946), .W4TO0(10), .W5TO0(-180), .W6TO0(-750), .W7TO0(-765), .W8TO0(916), .W9TO0(973), .W10TO0(779), .W11TO0(-737), .W12TO0(191), .W13TO0(-445), .W14TO0(311), .W15TO0(-969), .W16TO0(-172), .W17TO0(-606), .W18TO0(-19), .W19TO0(73), .W20TO0(669), .W21TO0(-147), .W22TO0(865), .W23TO0(-845), .W24TO0(-158), .W25TO0(837), .W26TO0(-713), .W27TO0(-402), .W28TO0(-158), .W29TO0(40), .W30TO0(-371), .W31TO0(577), .W32TO0(-85), .W33TO0(-501), .W34TO0(-220), .W35TO0(545), .W36TO0(-482), .W37TO0(-271), .W38TO0(-342), .W39TO0(-640), .W40TO0(767), .W41TO0(-506), .W42TO0(-804), .W43TO0(216), .W44TO0(992), .W45TO0(274), .W46TO0(551), .W47TO0(564), .W48TO0(-579), .W49TO0(-631), .W50TO0(141), .W51TO0(-562), .W52TO0(851), .W53TO0(208), .W54TO0(112), .W55TO0(-139), .W56TO0(-533), .W57TO0(304), .W58TO0(957), .W59TO0(220), .W60TO0(952), .W61TO0(-94), .W62TO0(-155), .W63TO0(20)) layer1(.clk(clk), .rst(rst), .in0(con0[0]), .in1(con0[1]), .in2(con0[2]), .in3(con0[3]), .in4(con0[4]), .in5(con0[5]), .in6(con0[6]), .in7(con0[7]), .in8(con0[8]), .in9(con0[9]), .in10(con0[10]), .in11(con0[11]), .in12(con0[12]), .in13(con0[13]), .in14(con0[14]), .in15(con0[15]), .in16(con0[16]), .in17(con0[17]), .in18(con0[18]), .in19(con0[19]), .in20(con0[20]), .in21(con0[21]), .in22(con0[22]), .in23(con0[23]), .in24(con0[24]), .in25(con0[25]), .in26(con0[26]), .in27(con0[27]), .in28(con0[28]), .in29(con0[29]), .in30(con0[30]), .in31(con0[31]), .in32(con0[32]), .in33(con0[33]), .in34(con0[34]), .in35(con0[35]), .in36(con0[36]), .in37(con0[37]), .in38(con0[38]), .in39(con0[39]), .in40(con0[40]), .in41(con0[41]), .in42(con0[42]), .in43(con0[43]), .in44(con0[44]), .in45(con0[45]), .in46(con0[46]), .in47(con0[47]), .in48(con0[48]), .in49(con0[49]), .in50(con0[50]), .in51(con0[51]), .in52(con0[52]), .in53(con0[53]), .in54(con0[54]), .in55(con0[55]), .in56(con0[56]), .in57(con0[57]), .in58(con0[58]), .in59(con0[59]), .in60(con0[60]), .in61(con0[61]), .in62(con0[62]), .in63(con0[63]), .out0(out0));

endmodule

`define assert_close(expected, got, eps) \
if ((expected > got && expected > got + eps) || (expected < got && expected + eps < got)) begin \
    $display("TEST FAILED in %m: got %d, expected %d", got, expected); \
end

module example_tb;
logic clk;
logic rst;

reg signed [15:0] net_in0, net_in1, net_in2, net_in3, net_in4, net_in5, net_in6, net_in7, net_in8, net_in9, net_in10, net_in11, net_in12, net_in13, net_in14, net_in15, net_in16, net_in17, net_in18, net_in19, net_in20, net_in21, net_in22, net_in23, net_in24, net_in25, net_in26, net_in27, net_in28, net_in29, net_in30, net_in31, net_in32, net_in33, net_in34, net_in35, net_in36, net_in37, net_in38, net_in39, net_in40, net_in41, net_in42, net_in43, net_in44, net_in45, net_in46, net_in47, net_in48, net_in49, net_in50, net_in51, net_in52, net_in53, net_in54, net_in55, net_in56, net_in57, net_in58, net_in59, net_in60, net_in61, net_in62, net_in63, net_in64;

wire signed [15:0] net_out0;

network net(.clk(clk), .rst(rst), .in0(net_in0), .in1(net_in1), .in2(net_in2), .in3(net_in3), .in4(net_in4), .in5(net_in5), .in6(net_in6), .in7(net_in7), .in8(net_in8), .in9(net_in9), .in10(net_in10), .in11(net_in11), .in12(net_in12), .in13(net_in13), .in14(net_in14), .in15(net_in15), .in16(net_in16), .in17(net_in17), .in18(net_in18), .in19(net_in19), .in20(net_in20), .in21(net_in21), .in22(net_in22), .in23(net_in23), .in24(net_in24), .in25(net_in25), .in26(net_in26), .in27(net_in27), .in28(net_in28), .in29(net_in29), .in30(net_in30), .in31(net_in31), .in32(net_in32), .in33(net_in33), .in34(net_in34), .in35(net_in35), .in36(net_in36), .in37(net_in37), .in38(net_in38), .in39(net_in39), .in40(net_in40), .in41(net_in41), .in42(net_in42), .in43(net_in43), .in44(net_in44), .in45(net_in45), .in46(net_in46), .in47(net_in47), .in48(net_in48), .in49(net_in49), .in50(net_in50), .in51(net_in51), .in52(net_in52), .in53(net_in53), .in54(net_in54), .in55(net_in55), .in56(net_in56), .in57(net_in57), .in58(net_in58), .in59(net_in59), .in60(net_in60), .in61(net_in61), .in62(net_in62), .in63(net_in63), .in64(net_in64), .out0(net_out0));

task test;
input signed [15:0] in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, out0;
begin
    net_in0 <= in0;
    net_in1 <= in1;
    net_in2 <= in2;
    net_in3 <= in3;
    net_in4 <= in4;
    net_in5 <= in5;
    net_in6 <= in6;
    net_in7 <= in7;
    net_in8 <= in8;
    net_in9 <= in9;
    net_in10 <= in10;
    net_in11 <= in11;
    net_in12 <= in12;
    net_in13 <= in13;
    net_in14 <= in14;
    net_in15 <= in15;
    net_in16 <= in16;
    net_in17 <= in17;
    net_in18 <= in18;
    net_in19 <= in19;
    net_in20 <= in20;
    net_in21 <= in21;
    net_in22 <= in22;
    net_in23 <= in23;
    net_in24 <= in24;
    net_in25 <= in25;
    net_in26 <= in26;
    net_in27 <= in27;
    net_in28 <= in28;
    net_in29 <= in29;
    net_in30 <= in30;
    net_in31 <= in31;
    net_in32 <= in32;
    net_in33 <= in33;
    net_in34 <= in34;
    net_in35 <= in35;
    net_in36 <= in36;
    net_in37 <= in37;
    net_in38 <= in38;
    net_in39 <= in39;
    net_in40 <= in40;
    net_in41 <= in41;
    net_in42 <= in42;
    net_in43 <= in43;
    net_in44 <= in44;
    net_in45 <= in45;
    net_in46 <= in46;
    net_in47 <= in47;
    net_in48 <= in48;
    net_in49 <= in49;
    net_in50 <= in50;
    net_in51 <= in51;
    net_in52 <= in52;
    net_in53 <= in53;
    net_in54 <= in54;
    net_in55 <= in55;
    net_in56 <= in56;
    net_in57 <= in57;
    net_in58 <= in58;
    net_in59 <= in59;
    net_in60 <= in60;
    net_in61 <= in61;
    net_in62 <= in62;
    net_in63 <= in63;
    net_in64 <= in64;
    #10000ns
    `assert_close(out0, net_out0, 10);
end
endtask

initial
begin
    $dumpfile("waves.vcd");
    $dumpvars;
    test(0, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 0, 1000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 0, 1000, 1000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 215);
    $display("Test0 completed");
    test(1000, 0, 0, 1000, 1000, 1000, 0, 0, 0, 0, 0, 0, 0, 1000, 0, 0, 1000, 0, 1000, 0, 0, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 0, 0, 0, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 160);
    $display("Test1 completed");
    test(0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 0, 0, 0, 1000, 1000, 627);
    $display("Test2 completed");
    test(0, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 0, 1000, 1000, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 0, 0, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 0, 1000, 0, 0, 59);
    $display("Test3 completed");
    test(1000, 0, 0, 0, 1000, 0, 0, 1000, 0, 0, 0, 1000, 0, 1000, 0, 1000, 0, 1000, 0, 0, 1000, 1000, 0, 0, 1000, 1000, 0, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 0, 0, 57);
    $display("Test4 completed");
    test(0, 0, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 0, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 0, 74);
    $display("Test5 completed");
    test(0, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 1000, 1000, 0, 597);
    $display("Test6 completed");
    test(1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 0, 0, 0, 1000, 0, 0, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 120);
    $display("Test7 completed");
    test(1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 0, 0, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 0, 1000, 1000, 0, 0, 0, 0, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 0, 131);
    $display("Test8 completed");
    test(0, 0, 1000, 0, 0, 0, 0, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 1000, 0, 0, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 67);
    $display("Test9 completed");
    test(1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 0, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 0, 1000, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 0, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 72);
    $display("Test10 completed");
    test(0, 1000, 0, 0, 0, 0, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 0, 0, 0, 1000, 0, 1000, 0, 1000, 0, 0, 1000, 0, 0, 0, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 0, 58);
    $display("Test11 completed");
    test(1000, 1000, 1000, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 0, 1000, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 293);
    $display("Test12 completed");
    test(1000, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 81);
    $display("Test13 completed");
    test(0, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 289);
    $display("Test14 completed");
    test(0, 0, 0, 0, 0, 1000, 0, 1000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 1000, 0, 0, 0, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 0, 1000, 1000, 0, 0, 0, 0, 1000, 0, 0, 0, 0, 1000, 0, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 76);
    $display("Test15 completed");
    test(0, 1000, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 0, 1000, 1000, 1000, 0, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 0, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 126);
    $display("Test16 completed");
    test(0, 1000, 0, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 0, 0, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 1000, 1000, 0, 1000, 81);
    $display("Test17 completed");
    test(0, 0, 0, 1000, 0, 1000, 0, 0, 0, 1000, 0, 0, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 0, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 290);
    $display("Test18 completed");
    test(1000, 0, 1000, 1000, 1000, 0, 0, 0, 0, 1000, 0, 0, 0, 0, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 0, 0, 0, 0, 1000, 0, 0, 1000, 1000, 0, 0, 0, 0, 1000, 0, 0, 1000, 1000, 115);
    $display("Test19 completed");
    test(1000, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 0, 0, 0, 0, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 0, 0, 0, 1000, 0, 1000, 0, 1000, 0, 0, 1000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1000, 1000, 0, 0, 136);
    $display("Test20 completed");
    test(0, 0, 1000, 0, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 0, 0, 0, 0, 0, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 1000, 0, 0, 0, 152);
    $display("Test21 completed");
    test(0, 0, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 0, 0, 0, 0, 0, 0, 1000, 324);
    $display("Test22 completed");
    test(1000, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 1000, 0, 0, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 0, 0, 1000, 1000, 0, 0, 0, 0, 1000, 0, 0, 0, 1000, 1000, 0, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 1000, 0, 1000, 0, 0, 0, 0, 522);
    $display("Test23 completed");
    test(1000, 1000, 1000, 0, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 1000, 1000, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 0, 0, 0, 0, 1000, 0, 1000, 0, 0, 664);
    $display("Test24 completed");
    test(0, 1000, 1000, 0, 0, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 0, 1000, 1000, 1000, 0, 1000, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 502);
    $display("Test25 completed");
    test(1000, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 0, 179);
    $display("Test26 completed");
    test(1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 1000, 1000, 0, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 0, 0, 0, 0, 1000, 0, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 0, 302);
    $display("Test27 completed");
    test(0, 1000, 0, 0, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 0, 0, 0, 1000, 0, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 142);
    $display("Test28 completed");
    test(0, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 1000, 0, 1000, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 466);
    $display("Test29 completed");
    test(0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 0, 78);
    $display("Test30 completed");
    test(1000, 0, 0, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 0, 0, 482);
    $display("Test31 completed");
    test(0, 1000, 0, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 163);
    $display("Test32 completed");
    test(0, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 0, 0, 1000, 1000, 0, 0, 0, 0, 0, 0, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 0, 0, 0, 1000, 0, 0, 1000, 1000, 218);
    $display("Test33 completed");
    test(0, 0, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 0, 1000, 0, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 1000, 0, 0, 0, 1000, 229);
    $display("Test34 completed");
    test(0, 0, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 1000, 0, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 0, 1000, 0, 1000, 332);
    $display("Test35 completed");
    test(0, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 1000, 0, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 0, 0, 1000, 0, 0, 0, 0, 0, 1000, 0, 0, 1000, 0, 0, 0, 0, 1000, 0, 0, 0, 0, 99);
    $display("Test36 completed");
    test(1000, 0, 0, 1000, 0, 0, 0, 0, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 164);
    $display("Test37 completed");
    test(1000, 1000, 0, 1000, 0, 0, 0, 0, 0, 1000, 0, 0, 0, 1000, 0, 1000, 0, 0, 0, 0, 0, 0, 0, 0, 1000, 1000, 0, 0, 0, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 0, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 108);
    $display("Test38 completed");
    test(1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 0, 1000, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 0, 0, 0, 1000, 1000, 0, 0, 0, 1000, 0, 0, 1000, 0, 0, 1000, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 254);
    $display("Test39 completed");
    test(1000, 1000, 1000, 0, 1000, 0, 1000, 0, 0, 1000, 0, 0, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 0, 1000, 0, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 1000, 0, 0, 0, 0, 0, 0, 1000, 1000, 0, 0, 1000, 1000, 359);
    $display("Test40 completed");
    test(0, 1000, 1000, 0, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 0, 0, 0, 0, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 0, 1000, 0, 0, 0, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 0, 0, 0, 0, 1000, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 1000, 1000, 70);
    $display("Test41 completed");
    test(1000, 0, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 0, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 0, 0, 0, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 130);
    $display("Test42 completed");
    test(0, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 0, 0, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 0, 0, 0, 1000, 0, 0, 1000, 0, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 0, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 0, 195);
    $display("Test43 completed");
    test(0, 1000, 0, 0, 0, 1000, 0, 1000, 0, 0, 1000, 0, 0, 1000, 0, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 0, 0, 0, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 348);
    $display("Test44 completed");
    test(1000, 0, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 0, 0, 0, 0, 1000, 0, 0, 1000, 156);
    $display("Test45 completed");
    test(1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 0, 0, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 0, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 9);
    $display("Test46 completed");
    test(0, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 0, 0, 1000, 0, 0, 0, 0, 1000, 0, 0, 0, 1000, 0, 0, 0, 0, 1000, 0, 1000, 0, 0, 0, 0, 0, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 0, 85);
    $display("Test47 completed");
    test(0, 1000, 1000, 0, 0, 0, 1000, 0, 1000, 0, 0, 0, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 0, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 0, 0, 0, 1000, 1000, 1000, 0, 0, 0, 0, 138);
    $display("Test48 completed");
    test(0, 0, 0, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 0, 1000, 0, 1000, 0, 0, 0, 0, 0, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 51);
    $display("Test49 completed");
    test(0, 0, 0, 0, 1000, 0, 1000, 1000, 0, 0, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 0, 0, 0, 1000, 0, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 1000, 0, 0, 78);
    $display("Test50 completed");
    test(1000, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 0, 0, 0, 0, 0, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 0, 0, 0, 0, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 157);
    $display("Test51 completed");
    test(0, 0, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 0, 1000, 0, 1000, 0, 1000, 0, 186);
    $display("Test52 completed");
    test(1000, 0, 0, 0, 0, 0, 0, 1000, 0, 0, 1000, 0, 0, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 0, 0, 0, 0, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 64);
    $display("Test53 completed");
    test(1000, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 0, 0, 0, 1000, 0, 0, 0, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 1000, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 188);
    $display("Test54 completed");
    test(1000, 1000, 0, 0, 0, 1000, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 0, 0, 0, 0, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 0, 0, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 0, 0, 1000, 0, 1000, 1000, 1000, 210);
    $display("Test55 completed");
    test(0, 1000, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 0, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 47);
    $display("Test56 completed");
    test(0, 1000, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 54);
    $display("Test57 completed");
    test(0, 1000, 1000, 0, 0, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 0, 0, 0, 1000, 0, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 1000, 0, 433);
    $display("Test58 completed");
    test(0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 0, 0, 0, 1000, 1000, 0, 0, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 0, 0, 1000, 0, 0, 0, 0, 1000, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 0, 0, 1000, 0, 1000, 1000, 0, 0, 0, 0, 0, 1000, 1000, 0, 1000, 778);
    $display("Test59 completed");
    test(1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 0, 1000, 1000, 0, 0, 0, 0, 331);
    $display("Test60 completed");
    test(0, 1000, 0, 1000, 0, 0, 0, 0, 1000, 0, 0, 1000, 0, 0, 1000, 0, 0, 1000, 0, 0, 0, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 0, 0, 0, 152);
    $display("Test61 completed");
    test(1000, 1000, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 0, 0, 0, 0, 0, 1000, 0, 1000, 0, 1000, 0, 0, 0, 0, 1000, 0, 0, 0, 1000, 0, 0, 1000, 0, 1000, 0, 0, 0, 1000, 1000, 0, 0, 0, 387);
    $display("Test62 completed");
    test(1000, 0, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 0, 0, 182);
    $display("Test63 completed");
    test(1000, 1000, 1000, 0, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 0, 0, 0, 1000, 1000, 239);
    $display("Test64 completed");
    test(0, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 0, 0, 1000, 268);
    $display("Test65 completed");
    test(1000, 0, 0, 1000, 0, 0, 0, 1000, 0, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 1000, 0, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 1000, 0, 1000, 0, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 683);
    $display("Test66 completed");
    test(1000, 0, 0, 1000, 0, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 1000, 1000, 0, 0, 1000, 0, 0, 0, 0, 1000, 0, 1000, 1000, 1000, 0, 0, 0, 0, 0, 1000, 0, 1000, 0, 0, 0, 0, 1000, 0, 0, 1000, 0, 0, 1000, 0, 0, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 1000, 59);
    $display("Test67 completed");
    test(0, 0, 0, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 0, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 1000, 0, 1000, 0, 0, 0, 0, 0, 1000, 0, 1000, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 1000, 1000, 0, 1000, 1000, 1000, 114);
    $display("Test68 completed");
    test(1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 0, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 1000, 0, 0, 1000, 1000, 0, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 1000, 39);
    $display("Test69 completed");
    test(0, 0, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 0, 99);
    $display("Test70 completed");
    test(0, 1000, 0, 0, 0, 0, 0, 0, 0, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 0, 1000, 785);
    $display("Test71 completed");
    test(0, 1000, 0, 0, 1000, 1000, 1000, 0, 1000, 0, 1000, 0, 1000, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 0, 0, 0, 0, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 115);
    $display("Test72 completed");
    test(0, 0, 1000, 0, 0, 0, 0, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 143);
    $display("Test73 completed");
    test(0, 0, 0, 0, 1000, 0, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 0, 0, 0, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 0, 0, 1000, 0, 1000, 705);
    $display("Test74 completed");
    test(1000, 0, 1000, 0, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 179);
    $display("Test75 completed");
    test(1000, 0, 0, 0, 1000, 0, 1000, 0, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 0, 0, 0, 0, 0, 1000, 0, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 0, 0, 1000, 1000, 0, 0, 0, 1000, 0, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 196);
    $display("Test76 completed");
    test(0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 0, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 0, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1000, 0, 0, 1000, 0, 1000, 1000, 0, 0, 0, 0, 0, 228);
    $display("Test77 completed");
    test(1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 1000, 1000, 0, 1000, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 0, 0, 0, 0, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 0, 60);
    $display("Test78 completed");
    test(1000, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 0, 0, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 0, 73);
    $display("Test79 completed");
    test(1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 0, 0, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 0, 0, 0, 0, 1000, 0, 0, 0, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 510);
    $display("Test80 completed");
    test(0, 0, 1000, 0, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 0, 0, 1000, 0, 0, 0, 1000, 0, 1000, 1000, 0, 1000, 257);
    $display("Test81 completed");
    test(1000, 0, 1000, 1000, 1000, 0, 0, 0, 0, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 0, 0, 0, 0, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 41);
    $display("Test82 completed");
    test(0, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 0, 0, 0, 0, 1000, 0, 1000, 0, 0, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 1000, 248);
    $display("Test83 completed");
    test(0, 1000, 0, 0, 0, 0, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 0, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 0, 0, 0, 1000, 0, 1000, 0, 0, 0, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 0, 1000, 0, 0, 354);
    $display("Test84 completed");
    test(0, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 1000, 166);
    $display("Test85 completed");
    test(0, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 0, 0, 1000, 0, 0, 0, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 0, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 0, 1000, 80);
    $display("Test86 completed");
    test(1000, 0, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 0, 1000, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 0, 1000, 0, 0, 0, 1000, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 0, 0, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 0, 0, 1000, 271);
    $display("Test87 completed");
    test(0, 0, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 0, 0, 0, 0, 0, 0, 0, 1000, 0, 0, 0, 1000, 1000, 0, 0, 0, 1000, 0, 0, 1000, 0, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 0, 0, 211);
    $display("Test88 completed");
    test(0, 0, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 1000, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 0, 0, 0, 0, 1000, 0, 1000, 1000, 0, 0, 0, 0, 1000, 676);
    $display("Test89 completed");
    test(1000, 1000, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 0, 166);
    $display("Test90 completed");
    test(0, 0, 1000, 1000, 0, 0, 0, 0, 0, 0, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 61);
    $display("Test91 completed");
    test(0, 0, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 0, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 391);
    $display("Test92 completed");
    test(0, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 1000, 0, 0, 1000, 1000, 0, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 0, 1000, 0, 0, 0, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 0, 0, 1000, 1000, 1000, 0, 1000, 0, 0, 0, 0, 1000, 0, 0, 0, 1000, 0, 0, 1000, 60);
    $display("Test93 completed");
    test(1000, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 0, 0, 0, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 0, 1000, 0, 0, 0, 1000, 0, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 0, 72);
    $display("Test94 completed");
    test(1000, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 1000, 0, 0, 1000, 0, 0, 0, 1000, 1000, 0, 0, 0, 0, 1000, 0, 0, 1000, 0, 0, 0, 1000, 1000, 0, 0, 1000, 0, 1000, 1000, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 0, 102);
    $display("Test95 completed");
    test(0, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 1000, 0, 0, 0, 0, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 0, 0, 0, 0, 0, 1000, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 50);
    $display("Test96 completed");
    test(1000, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 0, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 0, 1000, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 0, 0, 0, 0, 0, 0, 1000, 0, 0, 1000, 74);
    $display("Test97 completed");
    test(1000, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 0, 0, 1000, 1000, 0, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 1000, 0, 1000, 0, 1000, 1000, 0, 0, 0, 1000, 0, 1000, 1000, 1000, 1000, 1000, 0, 1000, 0, 0, 1000, 1000, 0, 0, 0, 0, 0, 0, 1000, 1000, 1000, 0, 0, 1000, 0, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 31);
    $display("Test98 completed");
    test(0, 1000, 0, 1000, 0, 0, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 0, 1000, 1000, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 1000, 0, 1000, 1000, 0, 0, 1000, 1000, 0, 0, 1000, 0, 0, 1000, 1000, 0, 0, 0, 0, 0, 1000, 1000, 1000, 1000, 0, 0, 0, 0, 1000, 230);
    $display("Test99 completed");
    $display("SUCCESS!");
end
endmodule
