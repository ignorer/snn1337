module neuron64in(clk, rst, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, out);

parameter W0 = 0;
parameter W1 = 0;
parameter W2 = 0;
parameter W3 = 0;
parameter W4 = 0;
parameter W5 = 0;
parameter W6 = 0;
parameter W7 = 0;
parameter W8 = 0;
parameter W9 = 0;
parameter W10 = 0;
parameter W11 = 0;
parameter W12 = 0;
parameter W13 = 0;
parameter W14 = 0;
parameter W15 = 0;
parameter W16 = 0;
parameter W17 = 0;
parameter W18 = 0;
parameter W19 = 0;
parameter W20 = 0;
parameter W21 = 0;
parameter W22 = 0;
parameter W23 = 0;
parameter W24 = 0;
parameter W25 = 0;
parameter W26 = 0;
parameter W27 = 0;
parameter W28 = 0;
parameter W29 = 0;
parameter W30 = 0;
parameter W31 = 0;
parameter W32 = 0;
parameter W33 = 0;
parameter W34 = 0;
parameter W35 = 0;
parameter W36 = 0;
parameter W37 = 0;
parameter W38 = 0;
parameter W39 = 0;
parameter W40 = 0;
parameter W41 = 0;
parameter W42 = 0;
parameter W43 = 0;
parameter W44 = 0;
parameter W45 = 0;
parameter W46 = 0;
parameter W47 = 0;
parameter W48 = 0;
parameter W49 = 0;
parameter W50 = 0;
parameter W51 = 0;
parameter W52 = 0;
parameter W53 = 0;
parameter W54 = 0;
parameter W55 = 0;
parameter W56 = 0;
parameter W57 = 0;
parameter W58 = 0;
parameter W59 = 0;
parameter W60 = 0;
parameter W61 = 0;
parameter W62 = 0;
parameter W63 = 0;

input wire clk;
input wire rst;

input signed [15:0] in0;
input signed [15:0] in1;
input signed [15:0] in2;
input signed [15:0] in3;
input signed [15:0] in4;
input signed [15:0] in5;
input signed [15:0] in6;
input signed [15:0] in7;
input signed [15:0] in8;
input signed [15:0] in9;
input signed [15:0] in10;
input signed [15:0] in11;
input signed [15:0] in12;
input signed [15:0] in13;
input signed [15:0] in14;
input signed [15:0] in15;
input signed [15:0] in16;
input signed [15:0] in17;
input signed [15:0] in18;
input signed [15:0] in19;
input signed [15:0] in20;
input signed [15:0] in21;
input signed [15:0] in22;
input signed [15:0] in23;
input signed [15:0] in24;
input signed [15:0] in25;
input signed [15:0] in26;
input signed [15:0] in27;
input signed [15:0] in28;
input signed [15:0] in29;
input signed [15:0] in30;
input signed [15:0] in31;
input signed [15:0] in32;
input signed [15:0] in33;
input signed [15:0] in34;
input signed [15:0] in35;
input signed [15:0] in36;
input signed [15:0] in37;
input signed [15:0] in38;
input signed [15:0] in39;
input signed [15:0] in40;
input signed [15:0] in41;
input signed [15:0] in42;
input signed [15:0] in43;
input signed [15:0] in44;
input signed [15:0] in45;
input signed [15:0] in46;
input signed [15:0] in47;
input signed [15:0] in48;
input signed [15:0] in49;
input signed [15:0] in50;
input signed [15:0] in51;
input signed [15:0] in52;
input signed [15:0] in53;
input signed [15:0] in54;
input signed [15:0] in55;
input signed [15:0] in56;
input signed [15:0] in57;
input signed [15:0] in58;
input signed [15:0] in59;
input signed [15:0] in60;
input signed [15:0] in61;
input signed [15:0] in62;
input signed [15:0] in63;

output reg signed [15:0] out;

reg signed [31:0] x;
reg [31:0] abs_x;
reg [31:0] y;
always @* begin
    x = in0 * W0 / 1000 + in1 * W1 / 1000 + in2 * W2 / 1000 + in3 * W3 / 1000 + in4 * W4 / 1000 + in5 * W5 / 1000 + in6 * W6 / 1000 + in7 * W7 / 1000 + in8 * W8 / 1000 + in9 * W9 / 1000 + in10 * W10 / 1000 + in11 * W11 / 1000 + in12 * W12 / 1000 + in13 * W13 / 1000 + in14 * W14 / 1000 + in15 * W15 / 1000 + in16 * W16 / 1000 + in17 * W17 / 1000 + in18 * W18 / 1000 + in19 * W19 / 1000 + in20 * W20 / 1000 + in21 * W21 / 1000 + in22 * W22 / 1000 + in23 * W23 / 1000 + in24 * W24 / 1000 + in25 * W25 / 1000 + in26 * W26 / 1000 + in27 * W27 / 1000 + in28 * W28 / 1000 + in29 * W29 / 1000 + in30 * W30 / 1000 + in31 * W31 / 1000 + in32 * W32 / 1000 + in33 * W33 / 1000 + in34 * W34 / 1000 + in35 * W35 / 1000 + in36 * W36 / 1000 + in37 * W37 / 1000 + in38 * W38 / 1000 + in39 * W39 / 1000 + in40 * W40 / 1000 + in41 * W41 / 1000 + in42 * W42 / 1000 + in43 * W43 / 1000 + in44 * W44 / 1000 + in45 * W45 / 1000 + in46 * W46 / 1000 + in47 * W47 / 1000 + in48 * W48 / 1000 + in49 * W49 / 1000 + in50 * W50 / 1000 + in51 * W51 / 1000 + in52 * W52 / 1000 + in53 * W53 / 1000 + in54 * W54 / 1000 + in55 * W55 / 1000 + in56 * W56 / 1000 + in57 * W57 / 1000 + in58 * W58 / 1000 + in59 * W59 / 1000 + in60 * W60 / 1000 + in61 * W61 / 1000 + in62 * W62 / 1000 + in63 * W63 / 1000;
    abs_x = x < 0 ? -x : x;
    if (abs_x >= 5000) y = 1000;
    else if (abs_x >= 2375) y = 31 * abs_x / 1000 + 844;
    else if (abs_x >= 1000) y = 125 * abs_x / 1000 + 625;
    else if (abs_x >= 0) y = 250 * abs_x / 1000 + 500;
    out = y;
end

endmodule

module neuron100in(clk, rst, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85, in86, in87, in88, in89, in90, in91, in92, in93, in94, in95, in96, in97, in98, in99, out);

parameter W0 = 0;
parameter W1 = 0;
parameter W2 = 0;
parameter W3 = 0;
parameter W4 = 0;
parameter W5 = 0;
parameter W6 = 0;
parameter W7 = 0;
parameter W8 = 0;
parameter W9 = 0;
parameter W10 = 0;
parameter W11 = 0;
parameter W12 = 0;
parameter W13 = 0;
parameter W14 = 0;
parameter W15 = 0;
parameter W16 = 0;
parameter W17 = 0;
parameter W18 = 0;
parameter W19 = 0;
parameter W20 = 0;
parameter W21 = 0;
parameter W22 = 0;
parameter W23 = 0;
parameter W24 = 0;
parameter W25 = 0;
parameter W26 = 0;
parameter W27 = 0;
parameter W28 = 0;
parameter W29 = 0;
parameter W30 = 0;
parameter W31 = 0;
parameter W32 = 0;
parameter W33 = 0;
parameter W34 = 0;
parameter W35 = 0;
parameter W36 = 0;
parameter W37 = 0;
parameter W38 = 0;
parameter W39 = 0;
parameter W40 = 0;
parameter W41 = 0;
parameter W42 = 0;
parameter W43 = 0;
parameter W44 = 0;
parameter W45 = 0;
parameter W46 = 0;
parameter W47 = 0;
parameter W48 = 0;
parameter W49 = 0;
parameter W50 = 0;
parameter W51 = 0;
parameter W52 = 0;
parameter W53 = 0;
parameter W54 = 0;
parameter W55 = 0;
parameter W56 = 0;
parameter W57 = 0;
parameter W58 = 0;
parameter W59 = 0;
parameter W60 = 0;
parameter W61 = 0;
parameter W62 = 0;
parameter W63 = 0;
parameter W64 = 0;
parameter W65 = 0;
parameter W66 = 0;
parameter W67 = 0;
parameter W68 = 0;
parameter W69 = 0;
parameter W70 = 0;
parameter W71 = 0;
parameter W72 = 0;
parameter W73 = 0;
parameter W74 = 0;
parameter W75 = 0;
parameter W76 = 0;
parameter W77 = 0;
parameter W78 = 0;
parameter W79 = 0;
parameter W80 = 0;
parameter W81 = 0;
parameter W82 = 0;
parameter W83 = 0;
parameter W84 = 0;
parameter W85 = 0;
parameter W86 = 0;
parameter W87 = 0;
parameter W88 = 0;
parameter W89 = 0;
parameter W90 = 0;
parameter W91 = 0;
parameter W92 = 0;
parameter W93 = 0;
parameter W94 = 0;
parameter W95 = 0;
parameter W96 = 0;
parameter W97 = 0;
parameter W98 = 0;
parameter W99 = 0;

input wire clk;
input wire rst;

input signed [15:0] in0;
input signed [15:0] in1;
input signed [15:0] in2;
input signed [15:0] in3;
input signed [15:0] in4;
input signed [15:0] in5;
input signed [15:0] in6;
input signed [15:0] in7;
input signed [15:0] in8;
input signed [15:0] in9;
input signed [15:0] in10;
input signed [15:0] in11;
input signed [15:0] in12;
input signed [15:0] in13;
input signed [15:0] in14;
input signed [15:0] in15;
input signed [15:0] in16;
input signed [15:0] in17;
input signed [15:0] in18;
input signed [15:0] in19;
input signed [15:0] in20;
input signed [15:0] in21;
input signed [15:0] in22;
input signed [15:0] in23;
input signed [15:0] in24;
input signed [15:0] in25;
input signed [15:0] in26;
input signed [15:0] in27;
input signed [15:0] in28;
input signed [15:0] in29;
input signed [15:0] in30;
input signed [15:0] in31;
input signed [15:0] in32;
input signed [15:0] in33;
input signed [15:0] in34;
input signed [15:0] in35;
input signed [15:0] in36;
input signed [15:0] in37;
input signed [15:0] in38;
input signed [15:0] in39;
input signed [15:0] in40;
input signed [15:0] in41;
input signed [15:0] in42;
input signed [15:0] in43;
input signed [15:0] in44;
input signed [15:0] in45;
input signed [15:0] in46;
input signed [15:0] in47;
input signed [15:0] in48;
input signed [15:0] in49;
input signed [15:0] in50;
input signed [15:0] in51;
input signed [15:0] in52;
input signed [15:0] in53;
input signed [15:0] in54;
input signed [15:0] in55;
input signed [15:0] in56;
input signed [15:0] in57;
input signed [15:0] in58;
input signed [15:0] in59;
input signed [15:0] in60;
input signed [15:0] in61;
input signed [15:0] in62;
input signed [15:0] in63;
input signed [15:0] in64;
input signed [15:0] in65;
input signed [15:0] in66;
input signed [15:0] in67;
input signed [15:0] in68;
input signed [15:0] in69;
input signed [15:0] in70;
input signed [15:0] in71;
input signed [15:0] in72;
input signed [15:0] in73;
input signed [15:0] in74;
input signed [15:0] in75;
input signed [15:0] in76;
input signed [15:0] in77;
input signed [15:0] in78;
input signed [15:0] in79;
input signed [15:0] in80;
input signed [15:0] in81;
input signed [15:0] in82;
input signed [15:0] in83;
input signed [15:0] in84;
input signed [15:0] in85;
input signed [15:0] in86;
input signed [15:0] in87;
input signed [15:0] in88;
input signed [15:0] in89;
input signed [15:0] in90;
input signed [15:0] in91;
input signed [15:0] in92;
input signed [15:0] in93;
input signed [15:0] in94;
input signed [15:0] in95;
input signed [15:0] in96;
input signed [15:0] in97;
input signed [15:0] in98;
input signed [15:0] in99;

output reg signed [15:0] out;

reg signed [31:0] x;
reg [31:0] abs_x;
reg [31:0] y;
always @* begin
    x = in0 * W0 / 1000 + in1 * W1 / 1000 + in2 * W2 / 1000 + in3 * W3 / 1000 + in4 * W4 / 1000 + in5 * W5 / 1000 + in6 * W6 / 1000 + in7 * W7 / 1000 + in8 * W8 / 1000 + in9 * W9 / 1000 + in10 * W10 / 1000 + in11 * W11 / 1000 + in12 * W12 / 1000 + in13 * W13 / 1000 + in14 * W14 / 1000 + in15 * W15 / 1000 + in16 * W16 / 1000 + in17 * W17 / 1000 + in18 * W18 / 1000 + in19 * W19 / 1000 + in20 * W20 / 1000 + in21 * W21 / 1000 + in22 * W22 / 1000 + in23 * W23 / 1000 + in24 * W24 / 1000 + in25 * W25 / 1000 + in26 * W26 / 1000 + in27 * W27 / 1000 + in28 * W28 / 1000 + in29 * W29 / 1000 + in30 * W30 / 1000 + in31 * W31 / 1000 + in32 * W32 / 1000 + in33 * W33 / 1000 + in34 * W34 / 1000 + in35 * W35 / 1000 + in36 * W36 / 1000 + in37 * W37 / 1000 + in38 * W38 / 1000 + in39 * W39 / 1000 + in40 * W40 / 1000 + in41 * W41 / 1000 + in42 * W42 / 1000 + in43 * W43 / 1000 + in44 * W44 / 1000 + in45 * W45 / 1000 + in46 * W46 / 1000 + in47 * W47 / 1000 + in48 * W48 / 1000 + in49 * W49 / 1000 + in50 * W50 / 1000 + in51 * W51 / 1000 + in52 * W52 / 1000 + in53 * W53 / 1000 + in54 * W54 / 1000 + in55 * W55 / 1000 + in56 * W56 / 1000 + in57 * W57 / 1000 + in58 * W58 / 1000 + in59 * W59 / 1000 + in60 * W60 / 1000 + in61 * W61 / 1000 + in62 * W62 / 1000 + in63 * W63 / 1000 + in64 * W64 / 1000 + in65 * W65 / 1000 + in66 * W66 / 1000 + in67 * W67 / 1000 + in68 * W68 / 1000 + in69 * W69 / 1000 + in70 * W70 / 1000 + in71 * W71 / 1000 + in72 * W72 / 1000 + in73 * W73 / 1000 + in74 * W74 / 1000 + in75 * W75 / 1000 + in76 * W76 / 1000 + in77 * W77 / 1000 + in78 * W78 / 1000 + in79 * W79 / 1000 + in80 * W80 / 1000 + in81 * W81 / 1000 + in82 * W82 / 1000 + in83 * W83 / 1000 + in84 * W84 / 1000 + in85 * W85 / 1000 + in86 * W86 / 1000 + in87 * W87 / 1000 + in88 * W88 / 1000 + in89 * W89 / 1000 + in90 * W90 / 1000 + in91 * W91 / 1000 + in92 * W92 / 1000 + in93 * W93 / 1000 + in94 * W94 / 1000 + in95 * W95 / 1000 + in96 * W96 / 1000 + in97 * W97 / 1000 + in98 * W98 / 1000 + in99 * W99 / 1000;
    abs_x = x < 0 ? -x : x;
    if (abs_x >= 5000) y = 1000;
    else if (abs_x >= 2375) y = 31 * abs_x / 1000 + 844;
    else if (abs_x >= 1000) y = 125 * abs_x / 1000 + 625;
    else if (abs_x >= 0) y = 250 * abs_x / 1000 + 500;
    out = y;
end

endmodule

module layer64in100out(clk, rst, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, out0, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13, out14, out15, out16, out17, out18, out19, out20, out21, out22, out23, out24, out25, out26, out27, out28, out29, out30, out31, out32, out33, out34, out35, out36, out37, out38, out39, out40, out41, out42, out43, out44, out45, out46, out47, out48, out49, out50, out51, out52, out53, out54, out55, out56, out57, out58, out59, out60, out61, out62, out63, out64, out65, out66, out67, out68, out69, out70, out71, out72, out73, out74, out75, out76, out77, out78, out79, out80, out81, out82, out83, out84, out85, out86, out87, out88, out89, out90, out91, out92, out93, out94, out95, out96, out97, out98, out99);

parameter W0TO0 = 0;
parameter W0TO1 = 0;
parameter W0TO2 = 0;
parameter W0TO3 = 0;
parameter W0TO4 = 0;
parameter W0TO5 = 0;
parameter W0TO6 = 0;
parameter W0TO7 = 0;
parameter W0TO8 = 0;
parameter W0TO9 = 0;
parameter W0TO10 = 0;
parameter W0TO11 = 0;
parameter W0TO12 = 0;
parameter W0TO13 = 0;
parameter W0TO14 = 0;
parameter W0TO15 = 0;
parameter W0TO16 = 0;
parameter W0TO17 = 0;
parameter W0TO18 = 0;
parameter W0TO19 = 0;
parameter W0TO20 = 0;
parameter W0TO21 = 0;
parameter W0TO22 = 0;
parameter W0TO23 = 0;
parameter W0TO24 = 0;
parameter W0TO25 = 0;
parameter W0TO26 = 0;
parameter W0TO27 = 0;
parameter W0TO28 = 0;
parameter W0TO29 = 0;
parameter W0TO30 = 0;
parameter W0TO31 = 0;
parameter W0TO32 = 0;
parameter W0TO33 = 0;
parameter W0TO34 = 0;
parameter W0TO35 = 0;
parameter W0TO36 = 0;
parameter W0TO37 = 0;
parameter W0TO38 = 0;
parameter W0TO39 = 0;
parameter W0TO40 = 0;
parameter W0TO41 = 0;
parameter W0TO42 = 0;
parameter W0TO43 = 0;
parameter W0TO44 = 0;
parameter W0TO45 = 0;
parameter W0TO46 = 0;
parameter W0TO47 = 0;
parameter W0TO48 = 0;
parameter W0TO49 = 0;
parameter W0TO50 = 0;
parameter W0TO51 = 0;
parameter W0TO52 = 0;
parameter W0TO53 = 0;
parameter W0TO54 = 0;
parameter W0TO55 = 0;
parameter W0TO56 = 0;
parameter W0TO57 = 0;
parameter W0TO58 = 0;
parameter W0TO59 = 0;
parameter W0TO60 = 0;
parameter W0TO61 = 0;
parameter W0TO62 = 0;
parameter W0TO63 = 0;
parameter W0TO64 = 0;
parameter W0TO65 = 0;
parameter W0TO66 = 0;
parameter W0TO67 = 0;
parameter W0TO68 = 0;
parameter W0TO69 = 0;
parameter W0TO70 = 0;
parameter W0TO71 = 0;
parameter W0TO72 = 0;
parameter W0TO73 = 0;
parameter W0TO74 = 0;
parameter W0TO75 = 0;
parameter W0TO76 = 0;
parameter W0TO77 = 0;
parameter W0TO78 = 0;
parameter W0TO79 = 0;
parameter W0TO80 = 0;
parameter W0TO81 = 0;
parameter W0TO82 = 0;
parameter W0TO83 = 0;
parameter W0TO84 = 0;
parameter W0TO85 = 0;
parameter W0TO86 = 0;
parameter W0TO87 = 0;
parameter W0TO88 = 0;
parameter W0TO89 = 0;
parameter W0TO90 = 0;
parameter W0TO91 = 0;
parameter W0TO92 = 0;
parameter W0TO93 = 0;
parameter W0TO94 = 0;
parameter W0TO95 = 0;
parameter W0TO96 = 0;
parameter W0TO97 = 0;
parameter W0TO98 = 0;
parameter W0TO99 = 0;
parameter W1TO0 = 0;
parameter W1TO1 = 0;
parameter W1TO2 = 0;
parameter W1TO3 = 0;
parameter W1TO4 = 0;
parameter W1TO5 = 0;
parameter W1TO6 = 0;
parameter W1TO7 = 0;
parameter W1TO8 = 0;
parameter W1TO9 = 0;
parameter W1TO10 = 0;
parameter W1TO11 = 0;
parameter W1TO12 = 0;
parameter W1TO13 = 0;
parameter W1TO14 = 0;
parameter W1TO15 = 0;
parameter W1TO16 = 0;
parameter W1TO17 = 0;
parameter W1TO18 = 0;
parameter W1TO19 = 0;
parameter W1TO20 = 0;
parameter W1TO21 = 0;
parameter W1TO22 = 0;
parameter W1TO23 = 0;
parameter W1TO24 = 0;
parameter W1TO25 = 0;
parameter W1TO26 = 0;
parameter W1TO27 = 0;
parameter W1TO28 = 0;
parameter W1TO29 = 0;
parameter W1TO30 = 0;
parameter W1TO31 = 0;
parameter W1TO32 = 0;
parameter W1TO33 = 0;
parameter W1TO34 = 0;
parameter W1TO35 = 0;
parameter W1TO36 = 0;
parameter W1TO37 = 0;
parameter W1TO38 = 0;
parameter W1TO39 = 0;
parameter W1TO40 = 0;
parameter W1TO41 = 0;
parameter W1TO42 = 0;
parameter W1TO43 = 0;
parameter W1TO44 = 0;
parameter W1TO45 = 0;
parameter W1TO46 = 0;
parameter W1TO47 = 0;
parameter W1TO48 = 0;
parameter W1TO49 = 0;
parameter W1TO50 = 0;
parameter W1TO51 = 0;
parameter W1TO52 = 0;
parameter W1TO53 = 0;
parameter W1TO54 = 0;
parameter W1TO55 = 0;
parameter W1TO56 = 0;
parameter W1TO57 = 0;
parameter W1TO58 = 0;
parameter W1TO59 = 0;
parameter W1TO60 = 0;
parameter W1TO61 = 0;
parameter W1TO62 = 0;
parameter W1TO63 = 0;
parameter W1TO64 = 0;
parameter W1TO65 = 0;
parameter W1TO66 = 0;
parameter W1TO67 = 0;
parameter W1TO68 = 0;
parameter W1TO69 = 0;
parameter W1TO70 = 0;
parameter W1TO71 = 0;
parameter W1TO72 = 0;
parameter W1TO73 = 0;
parameter W1TO74 = 0;
parameter W1TO75 = 0;
parameter W1TO76 = 0;
parameter W1TO77 = 0;
parameter W1TO78 = 0;
parameter W1TO79 = 0;
parameter W1TO80 = 0;
parameter W1TO81 = 0;
parameter W1TO82 = 0;
parameter W1TO83 = 0;
parameter W1TO84 = 0;
parameter W1TO85 = 0;
parameter W1TO86 = 0;
parameter W1TO87 = 0;
parameter W1TO88 = 0;
parameter W1TO89 = 0;
parameter W1TO90 = 0;
parameter W1TO91 = 0;
parameter W1TO92 = 0;
parameter W1TO93 = 0;
parameter W1TO94 = 0;
parameter W1TO95 = 0;
parameter W1TO96 = 0;
parameter W1TO97 = 0;
parameter W1TO98 = 0;
parameter W1TO99 = 0;
parameter W2TO0 = 0;
parameter W2TO1 = 0;
parameter W2TO2 = 0;
parameter W2TO3 = 0;
parameter W2TO4 = 0;
parameter W2TO5 = 0;
parameter W2TO6 = 0;
parameter W2TO7 = 0;
parameter W2TO8 = 0;
parameter W2TO9 = 0;
parameter W2TO10 = 0;
parameter W2TO11 = 0;
parameter W2TO12 = 0;
parameter W2TO13 = 0;
parameter W2TO14 = 0;
parameter W2TO15 = 0;
parameter W2TO16 = 0;
parameter W2TO17 = 0;
parameter W2TO18 = 0;
parameter W2TO19 = 0;
parameter W2TO20 = 0;
parameter W2TO21 = 0;
parameter W2TO22 = 0;
parameter W2TO23 = 0;
parameter W2TO24 = 0;
parameter W2TO25 = 0;
parameter W2TO26 = 0;
parameter W2TO27 = 0;
parameter W2TO28 = 0;
parameter W2TO29 = 0;
parameter W2TO30 = 0;
parameter W2TO31 = 0;
parameter W2TO32 = 0;
parameter W2TO33 = 0;
parameter W2TO34 = 0;
parameter W2TO35 = 0;
parameter W2TO36 = 0;
parameter W2TO37 = 0;
parameter W2TO38 = 0;
parameter W2TO39 = 0;
parameter W2TO40 = 0;
parameter W2TO41 = 0;
parameter W2TO42 = 0;
parameter W2TO43 = 0;
parameter W2TO44 = 0;
parameter W2TO45 = 0;
parameter W2TO46 = 0;
parameter W2TO47 = 0;
parameter W2TO48 = 0;
parameter W2TO49 = 0;
parameter W2TO50 = 0;
parameter W2TO51 = 0;
parameter W2TO52 = 0;
parameter W2TO53 = 0;
parameter W2TO54 = 0;
parameter W2TO55 = 0;
parameter W2TO56 = 0;
parameter W2TO57 = 0;
parameter W2TO58 = 0;
parameter W2TO59 = 0;
parameter W2TO60 = 0;
parameter W2TO61 = 0;
parameter W2TO62 = 0;
parameter W2TO63 = 0;
parameter W2TO64 = 0;
parameter W2TO65 = 0;
parameter W2TO66 = 0;
parameter W2TO67 = 0;
parameter W2TO68 = 0;
parameter W2TO69 = 0;
parameter W2TO70 = 0;
parameter W2TO71 = 0;
parameter W2TO72 = 0;
parameter W2TO73 = 0;
parameter W2TO74 = 0;
parameter W2TO75 = 0;
parameter W2TO76 = 0;
parameter W2TO77 = 0;
parameter W2TO78 = 0;
parameter W2TO79 = 0;
parameter W2TO80 = 0;
parameter W2TO81 = 0;
parameter W2TO82 = 0;
parameter W2TO83 = 0;
parameter W2TO84 = 0;
parameter W2TO85 = 0;
parameter W2TO86 = 0;
parameter W2TO87 = 0;
parameter W2TO88 = 0;
parameter W2TO89 = 0;
parameter W2TO90 = 0;
parameter W2TO91 = 0;
parameter W2TO92 = 0;
parameter W2TO93 = 0;
parameter W2TO94 = 0;
parameter W2TO95 = 0;
parameter W2TO96 = 0;
parameter W2TO97 = 0;
parameter W2TO98 = 0;
parameter W2TO99 = 0;
parameter W3TO0 = 0;
parameter W3TO1 = 0;
parameter W3TO2 = 0;
parameter W3TO3 = 0;
parameter W3TO4 = 0;
parameter W3TO5 = 0;
parameter W3TO6 = 0;
parameter W3TO7 = 0;
parameter W3TO8 = 0;
parameter W3TO9 = 0;
parameter W3TO10 = 0;
parameter W3TO11 = 0;
parameter W3TO12 = 0;
parameter W3TO13 = 0;
parameter W3TO14 = 0;
parameter W3TO15 = 0;
parameter W3TO16 = 0;
parameter W3TO17 = 0;
parameter W3TO18 = 0;
parameter W3TO19 = 0;
parameter W3TO20 = 0;
parameter W3TO21 = 0;
parameter W3TO22 = 0;
parameter W3TO23 = 0;
parameter W3TO24 = 0;
parameter W3TO25 = 0;
parameter W3TO26 = 0;
parameter W3TO27 = 0;
parameter W3TO28 = 0;
parameter W3TO29 = 0;
parameter W3TO30 = 0;
parameter W3TO31 = 0;
parameter W3TO32 = 0;
parameter W3TO33 = 0;
parameter W3TO34 = 0;
parameter W3TO35 = 0;
parameter W3TO36 = 0;
parameter W3TO37 = 0;
parameter W3TO38 = 0;
parameter W3TO39 = 0;
parameter W3TO40 = 0;
parameter W3TO41 = 0;
parameter W3TO42 = 0;
parameter W3TO43 = 0;
parameter W3TO44 = 0;
parameter W3TO45 = 0;
parameter W3TO46 = 0;
parameter W3TO47 = 0;
parameter W3TO48 = 0;
parameter W3TO49 = 0;
parameter W3TO50 = 0;
parameter W3TO51 = 0;
parameter W3TO52 = 0;
parameter W3TO53 = 0;
parameter W3TO54 = 0;
parameter W3TO55 = 0;
parameter W3TO56 = 0;
parameter W3TO57 = 0;
parameter W3TO58 = 0;
parameter W3TO59 = 0;
parameter W3TO60 = 0;
parameter W3TO61 = 0;
parameter W3TO62 = 0;
parameter W3TO63 = 0;
parameter W3TO64 = 0;
parameter W3TO65 = 0;
parameter W3TO66 = 0;
parameter W3TO67 = 0;
parameter W3TO68 = 0;
parameter W3TO69 = 0;
parameter W3TO70 = 0;
parameter W3TO71 = 0;
parameter W3TO72 = 0;
parameter W3TO73 = 0;
parameter W3TO74 = 0;
parameter W3TO75 = 0;
parameter W3TO76 = 0;
parameter W3TO77 = 0;
parameter W3TO78 = 0;
parameter W3TO79 = 0;
parameter W3TO80 = 0;
parameter W3TO81 = 0;
parameter W3TO82 = 0;
parameter W3TO83 = 0;
parameter W3TO84 = 0;
parameter W3TO85 = 0;
parameter W3TO86 = 0;
parameter W3TO87 = 0;
parameter W3TO88 = 0;
parameter W3TO89 = 0;
parameter W3TO90 = 0;
parameter W3TO91 = 0;
parameter W3TO92 = 0;
parameter W3TO93 = 0;
parameter W3TO94 = 0;
parameter W3TO95 = 0;
parameter W3TO96 = 0;
parameter W3TO97 = 0;
parameter W3TO98 = 0;
parameter W3TO99 = 0;
parameter W4TO0 = 0;
parameter W4TO1 = 0;
parameter W4TO2 = 0;
parameter W4TO3 = 0;
parameter W4TO4 = 0;
parameter W4TO5 = 0;
parameter W4TO6 = 0;
parameter W4TO7 = 0;
parameter W4TO8 = 0;
parameter W4TO9 = 0;
parameter W4TO10 = 0;
parameter W4TO11 = 0;
parameter W4TO12 = 0;
parameter W4TO13 = 0;
parameter W4TO14 = 0;
parameter W4TO15 = 0;
parameter W4TO16 = 0;
parameter W4TO17 = 0;
parameter W4TO18 = 0;
parameter W4TO19 = 0;
parameter W4TO20 = 0;
parameter W4TO21 = 0;
parameter W4TO22 = 0;
parameter W4TO23 = 0;
parameter W4TO24 = 0;
parameter W4TO25 = 0;
parameter W4TO26 = 0;
parameter W4TO27 = 0;
parameter W4TO28 = 0;
parameter W4TO29 = 0;
parameter W4TO30 = 0;
parameter W4TO31 = 0;
parameter W4TO32 = 0;
parameter W4TO33 = 0;
parameter W4TO34 = 0;
parameter W4TO35 = 0;
parameter W4TO36 = 0;
parameter W4TO37 = 0;
parameter W4TO38 = 0;
parameter W4TO39 = 0;
parameter W4TO40 = 0;
parameter W4TO41 = 0;
parameter W4TO42 = 0;
parameter W4TO43 = 0;
parameter W4TO44 = 0;
parameter W4TO45 = 0;
parameter W4TO46 = 0;
parameter W4TO47 = 0;
parameter W4TO48 = 0;
parameter W4TO49 = 0;
parameter W4TO50 = 0;
parameter W4TO51 = 0;
parameter W4TO52 = 0;
parameter W4TO53 = 0;
parameter W4TO54 = 0;
parameter W4TO55 = 0;
parameter W4TO56 = 0;
parameter W4TO57 = 0;
parameter W4TO58 = 0;
parameter W4TO59 = 0;
parameter W4TO60 = 0;
parameter W4TO61 = 0;
parameter W4TO62 = 0;
parameter W4TO63 = 0;
parameter W4TO64 = 0;
parameter W4TO65 = 0;
parameter W4TO66 = 0;
parameter W4TO67 = 0;
parameter W4TO68 = 0;
parameter W4TO69 = 0;
parameter W4TO70 = 0;
parameter W4TO71 = 0;
parameter W4TO72 = 0;
parameter W4TO73 = 0;
parameter W4TO74 = 0;
parameter W4TO75 = 0;
parameter W4TO76 = 0;
parameter W4TO77 = 0;
parameter W4TO78 = 0;
parameter W4TO79 = 0;
parameter W4TO80 = 0;
parameter W4TO81 = 0;
parameter W4TO82 = 0;
parameter W4TO83 = 0;
parameter W4TO84 = 0;
parameter W4TO85 = 0;
parameter W4TO86 = 0;
parameter W4TO87 = 0;
parameter W4TO88 = 0;
parameter W4TO89 = 0;
parameter W4TO90 = 0;
parameter W4TO91 = 0;
parameter W4TO92 = 0;
parameter W4TO93 = 0;
parameter W4TO94 = 0;
parameter W4TO95 = 0;
parameter W4TO96 = 0;
parameter W4TO97 = 0;
parameter W4TO98 = 0;
parameter W4TO99 = 0;
parameter W5TO0 = 0;
parameter W5TO1 = 0;
parameter W5TO2 = 0;
parameter W5TO3 = 0;
parameter W5TO4 = 0;
parameter W5TO5 = 0;
parameter W5TO6 = 0;
parameter W5TO7 = 0;
parameter W5TO8 = 0;
parameter W5TO9 = 0;
parameter W5TO10 = 0;
parameter W5TO11 = 0;
parameter W5TO12 = 0;
parameter W5TO13 = 0;
parameter W5TO14 = 0;
parameter W5TO15 = 0;
parameter W5TO16 = 0;
parameter W5TO17 = 0;
parameter W5TO18 = 0;
parameter W5TO19 = 0;
parameter W5TO20 = 0;
parameter W5TO21 = 0;
parameter W5TO22 = 0;
parameter W5TO23 = 0;
parameter W5TO24 = 0;
parameter W5TO25 = 0;
parameter W5TO26 = 0;
parameter W5TO27 = 0;
parameter W5TO28 = 0;
parameter W5TO29 = 0;
parameter W5TO30 = 0;
parameter W5TO31 = 0;
parameter W5TO32 = 0;
parameter W5TO33 = 0;
parameter W5TO34 = 0;
parameter W5TO35 = 0;
parameter W5TO36 = 0;
parameter W5TO37 = 0;
parameter W5TO38 = 0;
parameter W5TO39 = 0;
parameter W5TO40 = 0;
parameter W5TO41 = 0;
parameter W5TO42 = 0;
parameter W5TO43 = 0;
parameter W5TO44 = 0;
parameter W5TO45 = 0;
parameter W5TO46 = 0;
parameter W5TO47 = 0;
parameter W5TO48 = 0;
parameter W5TO49 = 0;
parameter W5TO50 = 0;
parameter W5TO51 = 0;
parameter W5TO52 = 0;
parameter W5TO53 = 0;
parameter W5TO54 = 0;
parameter W5TO55 = 0;
parameter W5TO56 = 0;
parameter W5TO57 = 0;
parameter W5TO58 = 0;
parameter W5TO59 = 0;
parameter W5TO60 = 0;
parameter W5TO61 = 0;
parameter W5TO62 = 0;
parameter W5TO63 = 0;
parameter W5TO64 = 0;
parameter W5TO65 = 0;
parameter W5TO66 = 0;
parameter W5TO67 = 0;
parameter W5TO68 = 0;
parameter W5TO69 = 0;
parameter W5TO70 = 0;
parameter W5TO71 = 0;
parameter W5TO72 = 0;
parameter W5TO73 = 0;
parameter W5TO74 = 0;
parameter W5TO75 = 0;
parameter W5TO76 = 0;
parameter W5TO77 = 0;
parameter W5TO78 = 0;
parameter W5TO79 = 0;
parameter W5TO80 = 0;
parameter W5TO81 = 0;
parameter W5TO82 = 0;
parameter W5TO83 = 0;
parameter W5TO84 = 0;
parameter W5TO85 = 0;
parameter W5TO86 = 0;
parameter W5TO87 = 0;
parameter W5TO88 = 0;
parameter W5TO89 = 0;
parameter W5TO90 = 0;
parameter W5TO91 = 0;
parameter W5TO92 = 0;
parameter W5TO93 = 0;
parameter W5TO94 = 0;
parameter W5TO95 = 0;
parameter W5TO96 = 0;
parameter W5TO97 = 0;
parameter W5TO98 = 0;
parameter W5TO99 = 0;
parameter W6TO0 = 0;
parameter W6TO1 = 0;
parameter W6TO2 = 0;
parameter W6TO3 = 0;
parameter W6TO4 = 0;
parameter W6TO5 = 0;
parameter W6TO6 = 0;
parameter W6TO7 = 0;
parameter W6TO8 = 0;
parameter W6TO9 = 0;
parameter W6TO10 = 0;
parameter W6TO11 = 0;
parameter W6TO12 = 0;
parameter W6TO13 = 0;
parameter W6TO14 = 0;
parameter W6TO15 = 0;
parameter W6TO16 = 0;
parameter W6TO17 = 0;
parameter W6TO18 = 0;
parameter W6TO19 = 0;
parameter W6TO20 = 0;
parameter W6TO21 = 0;
parameter W6TO22 = 0;
parameter W6TO23 = 0;
parameter W6TO24 = 0;
parameter W6TO25 = 0;
parameter W6TO26 = 0;
parameter W6TO27 = 0;
parameter W6TO28 = 0;
parameter W6TO29 = 0;
parameter W6TO30 = 0;
parameter W6TO31 = 0;
parameter W6TO32 = 0;
parameter W6TO33 = 0;
parameter W6TO34 = 0;
parameter W6TO35 = 0;
parameter W6TO36 = 0;
parameter W6TO37 = 0;
parameter W6TO38 = 0;
parameter W6TO39 = 0;
parameter W6TO40 = 0;
parameter W6TO41 = 0;
parameter W6TO42 = 0;
parameter W6TO43 = 0;
parameter W6TO44 = 0;
parameter W6TO45 = 0;
parameter W6TO46 = 0;
parameter W6TO47 = 0;
parameter W6TO48 = 0;
parameter W6TO49 = 0;
parameter W6TO50 = 0;
parameter W6TO51 = 0;
parameter W6TO52 = 0;
parameter W6TO53 = 0;
parameter W6TO54 = 0;
parameter W6TO55 = 0;
parameter W6TO56 = 0;
parameter W6TO57 = 0;
parameter W6TO58 = 0;
parameter W6TO59 = 0;
parameter W6TO60 = 0;
parameter W6TO61 = 0;
parameter W6TO62 = 0;
parameter W6TO63 = 0;
parameter W6TO64 = 0;
parameter W6TO65 = 0;
parameter W6TO66 = 0;
parameter W6TO67 = 0;
parameter W6TO68 = 0;
parameter W6TO69 = 0;
parameter W6TO70 = 0;
parameter W6TO71 = 0;
parameter W6TO72 = 0;
parameter W6TO73 = 0;
parameter W6TO74 = 0;
parameter W6TO75 = 0;
parameter W6TO76 = 0;
parameter W6TO77 = 0;
parameter W6TO78 = 0;
parameter W6TO79 = 0;
parameter W6TO80 = 0;
parameter W6TO81 = 0;
parameter W6TO82 = 0;
parameter W6TO83 = 0;
parameter W6TO84 = 0;
parameter W6TO85 = 0;
parameter W6TO86 = 0;
parameter W6TO87 = 0;
parameter W6TO88 = 0;
parameter W6TO89 = 0;
parameter W6TO90 = 0;
parameter W6TO91 = 0;
parameter W6TO92 = 0;
parameter W6TO93 = 0;
parameter W6TO94 = 0;
parameter W6TO95 = 0;
parameter W6TO96 = 0;
parameter W6TO97 = 0;
parameter W6TO98 = 0;
parameter W6TO99 = 0;
parameter W7TO0 = 0;
parameter W7TO1 = 0;
parameter W7TO2 = 0;
parameter W7TO3 = 0;
parameter W7TO4 = 0;
parameter W7TO5 = 0;
parameter W7TO6 = 0;
parameter W7TO7 = 0;
parameter W7TO8 = 0;
parameter W7TO9 = 0;
parameter W7TO10 = 0;
parameter W7TO11 = 0;
parameter W7TO12 = 0;
parameter W7TO13 = 0;
parameter W7TO14 = 0;
parameter W7TO15 = 0;
parameter W7TO16 = 0;
parameter W7TO17 = 0;
parameter W7TO18 = 0;
parameter W7TO19 = 0;
parameter W7TO20 = 0;
parameter W7TO21 = 0;
parameter W7TO22 = 0;
parameter W7TO23 = 0;
parameter W7TO24 = 0;
parameter W7TO25 = 0;
parameter W7TO26 = 0;
parameter W7TO27 = 0;
parameter W7TO28 = 0;
parameter W7TO29 = 0;
parameter W7TO30 = 0;
parameter W7TO31 = 0;
parameter W7TO32 = 0;
parameter W7TO33 = 0;
parameter W7TO34 = 0;
parameter W7TO35 = 0;
parameter W7TO36 = 0;
parameter W7TO37 = 0;
parameter W7TO38 = 0;
parameter W7TO39 = 0;
parameter W7TO40 = 0;
parameter W7TO41 = 0;
parameter W7TO42 = 0;
parameter W7TO43 = 0;
parameter W7TO44 = 0;
parameter W7TO45 = 0;
parameter W7TO46 = 0;
parameter W7TO47 = 0;
parameter W7TO48 = 0;
parameter W7TO49 = 0;
parameter W7TO50 = 0;
parameter W7TO51 = 0;
parameter W7TO52 = 0;
parameter W7TO53 = 0;
parameter W7TO54 = 0;
parameter W7TO55 = 0;
parameter W7TO56 = 0;
parameter W7TO57 = 0;
parameter W7TO58 = 0;
parameter W7TO59 = 0;
parameter W7TO60 = 0;
parameter W7TO61 = 0;
parameter W7TO62 = 0;
parameter W7TO63 = 0;
parameter W7TO64 = 0;
parameter W7TO65 = 0;
parameter W7TO66 = 0;
parameter W7TO67 = 0;
parameter W7TO68 = 0;
parameter W7TO69 = 0;
parameter W7TO70 = 0;
parameter W7TO71 = 0;
parameter W7TO72 = 0;
parameter W7TO73 = 0;
parameter W7TO74 = 0;
parameter W7TO75 = 0;
parameter W7TO76 = 0;
parameter W7TO77 = 0;
parameter W7TO78 = 0;
parameter W7TO79 = 0;
parameter W7TO80 = 0;
parameter W7TO81 = 0;
parameter W7TO82 = 0;
parameter W7TO83 = 0;
parameter W7TO84 = 0;
parameter W7TO85 = 0;
parameter W7TO86 = 0;
parameter W7TO87 = 0;
parameter W7TO88 = 0;
parameter W7TO89 = 0;
parameter W7TO90 = 0;
parameter W7TO91 = 0;
parameter W7TO92 = 0;
parameter W7TO93 = 0;
parameter W7TO94 = 0;
parameter W7TO95 = 0;
parameter W7TO96 = 0;
parameter W7TO97 = 0;
parameter W7TO98 = 0;
parameter W7TO99 = 0;
parameter W8TO0 = 0;
parameter W8TO1 = 0;
parameter W8TO2 = 0;
parameter W8TO3 = 0;
parameter W8TO4 = 0;
parameter W8TO5 = 0;
parameter W8TO6 = 0;
parameter W8TO7 = 0;
parameter W8TO8 = 0;
parameter W8TO9 = 0;
parameter W8TO10 = 0;
parameter W8TO11 = 0;
parameter W8TO12 = 0;
parameter W8TO13 = 0;
parameter W8TO14 = 0;
parameter W8TO15 = 0;
parameter W8TO16 = 0;
parameter W8TO17 = 0;
parameter W8TO18 = 0;
parameter W8TO19 = 0;
parameter W8TO20 = 0;
parameter W8TO21 = 0;
parameter W8TO22 = 0;
parameter W8TO23 = 0;
parameter W8TO24 = 0;
parameter W8TO25 = 0;
parameter W8TO26 = 0;
parameter W8TO27 = 0;
parameter W8TO28 = 0;
parameter W8TO29 = 0;
parameter W8TO30 = 0;
parameter W8TO31 = 0;
parameter W8TO32 = 0;
parameter W8TO33 = 0;
parameter W8TO34 = 0;
parameter W8TO35 = 0;
parameter W8TO36 = 0;
parameter W8TO37 = 0;
parameter W8TO38 = 0;
parameter W8TO39 = 0;
parameter W8TO40 = 0;
parameter W8TO41 = 0;
parameter W8TO42 = 0;
parameter W8TO43 = 0;
parameter W8TO44 = 0;
parameter W8TO45 = 0;
parameter W8TO46 = 0;
parameter W8TO47 = 0;
parameter W8TO48 = 0;
parameter W8TO49 = 0;
parameter W8TO50 = 0;
parameter W8TO51 = 0;
parameter W8TO52 = 0;
parameter W8TO53 = 0;
parameter W8TO54 = 0;
parameter W8TO55 = 0;
parameter W8TO56 = 0;
parameter W8TO57 = 0;
parameter W8TO58 = 0;
parameter W8TO59 = 0;
parameter W8TO60 = 0;
parameter W8TO61 = 0;
parameter W8TO62 = 0;
parameter W8TO63 = 0;
parameter W8TO64 = 0;
parameter W8TO65 = 0;
parameter W8TO66 = 0;
parameter W8TO67 = 0;
parameter W8TO68 = 0;
parameter W8TO69 = 0;
parameter W8TO70 = 0;
parameter W8TO71 = 0;
parameter W8TO72 = 0;
parameter W8TO73 = 0;
parameter W8TO74 = 0;
parameter W8TO75 = 0;
parameter W8TO76 = 0;
parameter W8TO77 = 0;
parameter W8TO78 = 0;
parameter W8TO79 = 0;
parameter W8TO80 = 0;
parameter W8TO81 = 0;
parameter W8TO82 = 0;
parameter W8TO83 = 0;
parameter W8TO84 = 0;
parameter W8TO85 = 0;
parameter W8TO86 = 0;
parameter W8TO87 = 0;
parameter W8TO88 = 0;
parameter W8TO89 = 0;
parameter W8TO90 = 0;
parameter W8TO91 = 0;
parameter W8TO92 = 0;
parameter W8TO93 = 0;
parameter W8TO94 = 0;
parameter W8TO95 = 0;
parameter W8TO96 = 0;
parameter W8TO97 = 0;
parameter W8TO98 = 0;
parameter W8TO99 = 0;
parameter W9TO0 = 0;
parameter W9TO1 = 0;
parameter W9TO2 = 0;
parameter W9TO3 = 0;
parameter W9TO4 = 0;
parameter W9TO5 = 0;
parameter W9TO6 = 0;
parameter W9TO7 = 0;
parameter W9TO8 = 0;
parameter W9TO9 = 0;
parameter W9TO10 = 0;
parameter W9TO11 = 0;
parameter W9TO12 = 0;
parameter W9TO13 = 0;
parameter W9TO14 = 0;
parameter W9TO15 = 0;
parameter W9TO16 = 0;
parameter W9TO17 = 0;
parameter W9TO18 = 0;
parameter W9TO19 = 0;
parameter W9TO20 = 0;
parameter W9TO21 = 0;
parameter W9TO22 = 0;
parameter W9TO23 = 0;
parameter W9TO24 = 0;
parameter W9TO25 = 0;
parameter W9TO26 = 0;
parameter W9TO27 = 0;
parameter W9TO28 = 0;
parameter W9TO29 = 0;
parameter W9TO30 = 0;
parameter W9TO31 = 0;
parameter W9TO32 = 0;
parameter W9TO33 = 0;
parameter W9TO34 = 0;
parameter W9TO35 = 0;
parameter W9TO36 = 0;
parameter W9TO37 = 0;
parameter W9TO38 = 0;
parameter W9TO39 = 0;
parameter W9TO40 = 0;
parameter W9TO41 = 0;
parameter W9TO42 = 0;
parameter W9TO43 = 0;
parameter W9TO44 = 0;
parameter W9TO45 = 0;
parameter W9TO46 = 0;
parameter W9TO47 = 0;
parameter W9TO48 = 0;
parameter W9TO49 = 0;
parameter W9TO50 = 0;
parameter W9TO51 = 0;
parameter W9TO52 = 0;
parameter W9TO53 = 0;
parameter W9TO54 = 0;
parameter W9TO55 = 0;
parameter W9TO56 = 0;
parameter W9TO57 = 0;
parameter W9TO58 = 0;
parameter W9TO59 = 0;
parameter W9TO60 = 0;
parameter W9TO61 = 0;
parameter W9TO62 = 0;
parameter W9TO63 = 0;
parameter W9TO64 = 0;
parameter W9TO65 = 0;
parameter W9TO66 = 0;
parameter W9TO67 = 0;
parameter W9TO68 = 0;
parameter W9TO69 = 0;
parameter W9TO70 = 0;
parameter W9TO71 = 0;
parameter W9TO72 = 0;
parameter W9TO73 = 0;
parameter W9TO74 = 0;
parameter W9TO75 = 0;
parameter W9TO76 = 0;
parameter W9TO77 = 0;
parameter W9TO78 = 0;
parameter W9TO79 = 0;
parameter W9TO80 = 0;
parameter W9TO81 = 0;
parameter W9TO82 = 0;
parameter W9TO83 = 0;
parameter W9TO84 = 0;
parameter W9TO85 = 0;
parameter W9TO86 = 0;
parameter W9TO87 = 0;
parameter W9TO88 = 0;
parameter W9TO89 = 0;
parameter W9TO90 = 0;
parameter W9TO91 = 0;
parameter W9TO92 = 0;
parameter W9TO93 = 0;
parameter W9TO94 = 0;
parameter W9TO95 = 0;
parameter W9TO96 = 0;
parameter W9TO97 = 0;
parameter W9TO98 = 0;
parameter W9TO99 = 0;
parameter W10TO0 = 0;
parameter W10TO1 = 0;
parameter W10TO2 = 0;
parameter W10TO3 = 0;
parameter W10TO4 = 0;
parameter W10TO5 = 0;
parameter W10TO6 = 0;
parameter W10TO7 = 0;
parameter W10TO8 = 0;
parameter W10TO9 = 0;
parameter W10TO10 = 0;
parameter W10TO11 = 0;
parameter W10TO12 = 0;
parameter W10TO13 = 0;
parameter W10TO14 = 0;
parameter W10TO15 = 0;
parameter W10TO16 = 0;
parameter W10TO17 = 0;
parameter W10TO18 = 0;
parameter W10TO19 = 0;
parameter W10TO20 = 0;
parameter W10TO21 = 0;
parameter W10TO22 = 0;
parameter W10TO23 = 0;
parameter W10TO24 = 0;
parameter W10TO25 = 0;
parameter W10TO26 = 0;
parameter W10TO27 = 0;
parameter W10TO28 = 0;
parameter W10TO29 = 0;
parameter W10TO30 = 0;
parameter W10TO31 = 0;
parameter W10TO32 = 0;
parameter W10TO33 = 0;
parameter W10TO34 = 0;
parameter W10TO35 = 0;
parameter W10TO36 = 0;
parameter W10TO37 = 0;
parameter W10TO38 = 0;
parameter W10TO39 = 0;
parameter W10TO40 = 0;
parameter W10TO41 = 0;
parameter W10TO42 = 0;
parameter W10TO43 = 0;
parameter W10TO44 = 0;
parameter W10TO45 = 0;
parameter W10TO46 = 0;
parameter W10TO47 = 0;
parameter W10TO48 = 0;
parameter W10TO49 = 0;
parameter W10TO50 = 0;
parameter W10TO51 = 0;
parameter W10TO52 = 0;
parameter W10TO53 = 0;
parameter W10TO54 = 0;
parameter W10TO55 = 0;
parameter W10TO56 = 0;
parameter W10TO57 = 0;
parameter W10TO58 = 0;
parameter W10TO59 = 0;
parameter W10TO60 = 0;
parameter W10TO61 = 0;
parameter W10TO62 = 0;
parameter W10TO63 = 0;
parameter W10TO64 = 0;
parameter W10TO65 = 0;
parameter W10TO66 = 0;
parameter W10TO67 = 0;
parameter W10TO68 = 0;
parameter W10TO69 = 0;
parameter W10TO70 = 0;
parameter W10TO71 = 0;
parameter W10TO72 = 0;
parameter W10TO73 = 0;
parameter W10TO74 = 0;
parameter W10TO75 = 0;
parameter W10TO76 = 0;
parameter W10TO77 = 0;
parameter W10TO78 = 0;
parameter W10TO79 = 0;
parameter W10TO80 = 0;
parameter W10TO81 = 0;
parameter W10TO82 = 0;
parameter W10TO83 = 0;
parameter W10TO84 = 0;
parameter W10TO85 = 0;
parameter W10TO86 = 0;
parameter W10TO87 = 0;
parameter W10TO88 = 0;
parameter W10TO89 = 0;
parameter W10TO90 = 0;
parameter W10TO91 = 0;
parameter W10TO92 = 0;
parameter W10TO93 = 0;
parameter W10TO94 = 0;
parameter W10TO95 = 0;
parameter W10TO96 = 0;
parameter W10TO97 = 0;
parameter W10TO98 = 0;
parameter W10TO99 = 0;
parameter W11TO0 = 0;
parameter W11TO1 = 0;
parameter W11TO2 = 0;
parameter W11TO3 = 0;
parameter W11TO4 = 0;
parameter W11TO5 = 0;
parameter W11TO6 = 0;
parameter W11TO7 = 0;
parameter W11TO8 = 0;
parameter W11TO9 = 0;
parameter W11TO10 = 0;
parameter W11TO11 = 0;
parameter W11TO12 = 0;
parameter W11TO13 = 0;
parameter W11TO14 = 0;
parameter W11TO15 = 0;
parameter W11TO16 = 0;
parameter W11TO17 = 0;
parameter W11TO18 = 0;
parameter W11TO19 = 0;
parameter W11TO20 = 0;
parameter W11TO21 = 0;
parameter W11TO22 = 0;
parameter W11TO23 = 0;
parameter W11TO24 = 0;
parameter W11TO25 = 0;
parameter W11TO26 = 0;
parameter W11TO27 = 0;
parameter W11TO28 = 0;
parameter W11TO29 = 0;
parameter W11TO30 = 0;
parameter W11TO31 = 0;
parameter W11TO32 = 0;
parameter W11TO33 = 0;
parameter W11TO34 = 0;
parameter W11TO35 = 0;
parameter W11TO36 = 0;
parameter W11TO37 = 0;
parameter W11TO38 = 0;
parameter W11TO39 = 0;
parameter W11TO40 = 0;
parameter W11TO41 = 0;
parameter W11TO42 = 0;
parameter W11TO43 = 0;
parameter W11TO44 = 0;
parameter W11TO45 = 0;
parameter W11TO46 = 0;
parameter W11TO47 = 0;
parameter W11TO48 = 0;
parameter W11TO49 = 0;
parameter W11TO50 = 0;
parameter W11TO51 = 0;
parameter W11TO52 = 0;
parameter W11TO53 = 0;
parameter W11TO54 = 0;
parameter W11TO55 = 0;
parameter W11TO56 = 0;
parameter W11TO57 = 0;
parameter W11TO58 = 0;
parameter W11TO59 = 0;
parameter W11TO60 = 0;
parameter W11TO61 = 0;
parameter W11TO62 = 0;
parameter W11TO63 = 0;
parameter W11TO64 = 0;
parameter W11TO65 = 0;
parameter W11TO66 = 0;
parameter W11TO67 = 0;
parameter W11TO68 = 0;
parameter W11TO69 = 0;
parameter W11TO70 = 0;
parameter W11TO71 = 0;
parameter W11TO72 = 0;
parameter W11TO73 = 0;
parameter W11TO74 = 0;
parameter W11TO75 = 0;
parameter W11TO76 = 0;
parameter W11TO77 = 0;
parameter W11TO78 = 0;
parameter W11TO79 = 0;
parameter W11TO80 = 0;
parameter W11TO81 = 0;
parameter W11TO82 = 0;
parameter W11TO83 = 0;
parameter W11TO84 = 0;
parameter W11TO85 = 0;
parameter W11TO86 = 0;
parameter W11TO87 = 0;
parameter W11TO88 = 0;
parameter W11TO89 = 0;
parameter W11TO90 = 0;
parameter W11TO91 = 0;
parameter W11TO92 = 0;
parameter W11TO93 = 0;
parameter W11TO94 = 0;
parameter W11TO95 = 0;
parameter W11TO96 = 0;
parameter W11TO97 = 0;
parameter W11TO98 = 0;
parameter W11TO99 = 0;
parameter W12TO0 = 0;
parameter W12TO1 = 0;
parameter W12TO2 = 0;
parameter W12TO3 = 0;
parameter W12TO4 = 0;
parameter W12TO5 = 0;
parameter W12TO6 = 0;
parameter W12TO7 = 0;
parameter W12TO8 = 0;
parameter W12TO9 = 0;
parameter W12TO10 = 0;
parameter W12TO11 = 0;
parameter W12TO12 = 0;
parameter W12TO13 = 0;
parameter W12TO14 = 0;
parameter W12TO15 = 0;
parameter W12TO16 = 0;
parameter W12TO17 = 0;
parameter W12TO18 = 0;
parameter W12TO19 = 0;
parameter W12TO20 = 0;
parameter W12TO21 = 0;
parameter W12TO22 = 0;
parameter W12TO23 = 0;
parameter W12TO24 = 0;
parameter W12TO25 = 0;
parameter W12TO26 = 0;
parameter W12TO27 = 0;
parameter W12TO28 = 0;
parameter W12TO29 = 0;
parameter W12TO30 = 0;
parameter W12TO31 = 0;
parameter W12TO32 = 0;
parameter W12TO33 = 0;
parameter W12TO34 = 0;
parameter W12TO35 = 0;
parameter W12TO36 = 0;
parameter W12TO37 = 0;
parameter W12TO38 = 0;
parameter W12TO39 = 0;
parameter W12TO40 = 0;
parameter W12TO41 = 0;
parameter W12TO42 = 0;
parameter W12TO43 = 0;
parameter W12TO44 = 0;
parameter W12TO45 = 0;
parameter W12TO46 = 0;
parameter W12TO47 = 0;
parameter W12TO48 = 0;
parameter W12TO49 = 0;
parameter W12TO50 = 0;
parameter W12TO51 = 0;
parameter W12TO52 = 0;
parameter W12TO53 = 0;
parameter W12TO54 = 0;
parameter W12TO55 = 0;
parameter W12TO56 = 0;
parameter W12TO57 = 0;
parameter W12TO58 = 0;
parameter W12TO59 = 0;
parameter W12TO60 = 0;
parameter W12TO61 = 0;
parameter W12TO62 = 0;
parameter W12TO63 = 0;
parameter W12TO64 = 0;
parameter W12TO65 = 0;
parameter W12TO66 = 0;
parameter W12TO67 = 0;
parameter W12TO68 = 0;
parameter W12TO69 = 0;
parameter W12TO70 = 0;
parameter W12TO71 = 0;
parameter W12TO72 = 0;
parameter W12TO73 = 0;
parameter W12TO74 = 0;
parameter W12TO75 = 0;
parameter W12TO76 = 0;
parameter W12TO77 = 0;
parameter W12TO78 = 0;
parameter W12TO79 = 0;
parameter W12TO80 = 0;
parameter W12TO81 = 0;
parameter W12TO82 = 0;
parameter W12TO83 = 0;
parameter W12TO84 = 0;
parameter W12TO85 = 0;
parameter W12TO86 = 0;
parameter W12TO87 = 0;
parameter W12TO88 = 0;
parameter W12TO89 = 0;
parameter W12TO90 = 0;
parameter W12TO91 = 0;
parameter W12TO92 = 0;
parameter W12TO93 = 0;
parameter W12TO94 = 0;
parameter W12TO95 = 0;
parameter W12TO96 = 0;
parameter W12TO97 = 0;
parameter W12TO98 = 0;
parameter W12TO99 = 0;
parameter W13TO0 = 0;
parameter W13TO1 = 0;
parameter W13TO2 = 0;
parameter W13TO3 = 0;
parameter W13TO4 = 0;
parameter W13TO5 = 0;
parameter W13TO6 = 0;
parameter W13TO7 = 0;
parameter W13TO8 = 0;
parameter W13TO9 = 0;
parameter W13TO10 = 0;
parameter W13TO11 = 0;
parameter W13TO12 = 0;
parameter W13TO13 = 0;
parameter W13TO14 = 0;
parameter W13TO15 = 0;
parameter W13TO16 = 0;
parameter W13TO17 = 0;
parameter W13TO18 = 0;
parameter W13TO19 = 0;
parameter W13TO20 = 0;
parameter W13TO21 = 0;
parameter W13TO22 = 0;
parameter W13TO23 = 0;
parameter W13TO24 = 0;
parameter W13TO25 = 0;
parameter W13TO26 = 0;
parameter W13TO27 = 0;
parameter W13TO28 = 0;
parameter W13TO29 = 0;
parameter W13TO30 = 0;
parameter W13TO31 = 0;
parameter W13TO32 = 0;
parameter W13TO33 = 0;
parameter W13TO34 = 0;
parameter W13TO35 = 0;
parameter W13TO36 = 0;
parameter W13TO37 = 0;
parameter W13TO38 = 0;
parameter W13TO39 = 0;
parameter W13TO40 = 0;
parameter W13TO41 = 0;
parameter W13TO42 = 0;
parameter W13TO43 = 0;
parameter W13TO44 = 0;
parameter W13TO45 = 0;
parameter W13TO46 = 0;
parameter W13TO47 = 0;
parameter W13TO48 = 0;
parameter W13TO49 = 0;
parameter W13TO50 = 0;
parameter W13TO51 = 0;
parameter W13TO52 = 0;
parameter W13TO53 = 0;
parameter W13TO54 = 0;
parameter W13TO55 = 0;
parameter W13TO56 = 0;
parameter W13TO57 = 0;
parameter W13TO58 = 0;
parameter W13TO59 = 0;
parameter W13TO60 = 0;
parameter W13TO61 = 0;
parameter W13TO62 = 0;
parameter W13TO63 = 0;
parameter W13TO64 = 0;
parameter W13TO65 = 0;
parameter W13TO66 = 0;
parameter W13TO67 = 0;
parameter W13TO68 = 0;
parameter W13TO69 = 0;
parameter W13TO70 = 0;
parameter W13TO71 = 0;
parameter W13TO72 = 0;
parameter W13TO73 = 0;
parameter W13TO74 = 0;
parameter W13TO75 = 0;
parameter W13TO76 = 0;
parameter W13TO77 = 0;
parameter W13TO78 = 0;
parameter W13TO79 = 0;
parameter W13TO80 = 0;
parameter W13TO81 = 0;
parameter W13TO82 = 0;
parameter W13TO83 = 0;
parameter W13TO84 = 0;
parameter W13TO85 = 0;
parameter W13TO86 = 0;
parameter W13TO87 = 0;
parameter W13TO88 = 0;
parameter W13TO89 = 0;
parameter W13TO90 = 0;
parameter W13TO91 = 0;
parameter W13TO92 = 0;
parameter W13TO93 = 0;
parameter W13TO94 = 0;
parameter W13TO95 = 0;
parameter W13TO96 = 0;
parameter W13TO97 = 0;
parameter W13TO98 = 0;
parameter W13TO99 = 0;
parameter W14TO0 = 0;
parameter W14TO1 = 0;
parameter W14TO2 = 0;
parameter W14TO3 = 0;
parameter W14TO4 = 0;
parameter W14TO5 = 0;
parameter W14TO6 = 0;
parameter W14TO7 = 0;
parameter W14TO8 = 0;
parameter W14TO9 = 0;
parameter W14TO10 = 0;
parameter W14TO11 = 0;
parameter W14TO12 = 0;
parameter W14TO13 = 0;
parameter W14TO14 = 0;
parameter W14TO15 = 0;
parameter W14TO16 = 0;
parameter W14TO17 = 0;
parameter W14TO18 = 0;
parameter W14TO19 = 0;
parameter W14TO20 = 0;
parameter W14TO21 = 0;
parameter W14TO22 = 0;
parameter W14TO23 = 0;
parameter W14TO24 = 0;
parameter W14TO25 = 0;
parameter W14TO26 = 0;
parameter W14TO27 = 0;
parameter W14TO28 = 0;
parameter W14TO29 = 0;
parameter W14TO30 = 0;
parameter W14TO31 = 0;
parameter W14TO32 = 0;
parameter W14TO33 = 0;
parameter W14TO34 = 0;
parameter W14TO35 = 0;
parameter W14TO36 = 0;
parameter W14TO37 = 0;
parameter W14TO38 = 0;
parameter W14TO39 = 0;
parameter W14TO40 = 0;
parameter W14TO41 = 0;
parameter W14TO42 = 0;
parameter W14TO43 = 0;
parameter W14TO44 = 0;
parameter W14TO45 = 0;
parameter W14TO46 = 0;
parameter W14TO47 = 0;
parameter W14TO48 = 0;
parameter W14TO49 = 0;
parameter W14TO50 = 0;
parameter W14TO51 = 0;
parameter W14TO52 = 0;
parameter W14TO53 = 0;
parameter W14TO54 = 0;
parameter W14TO55 = 0;
parameter W14TO56 = 0;
parameter W14TO57 = 0;
parameter W14TO58 = 0;
parameter W14TO59 = 0;
parameter W14TO60 = 0;
parameter W14TO61 = 0;
parameter W14TO62 = 0;
parameter W14TO63 = 0;
parameter W14TO64 = 0;
parameter W14TO65 = 0;
parameter W14TO66 = 0;
parameter W14TO67 = 0;
parameter W14TO68 = 0;
parameter W14TO69 = 0;
parameter W14TO70 = 0;
parameter W14TO71 = 0;
parameter W14TO72 = 0;
parameter W14TO73 = 0;
parameter W14TO74 = 0;
parameter W14TO75 = 0;
parameter W14TO76 = 0;
parameter W14TO77 = 0;
parameter W14TO78 = 0;
parameter W14TO79 = 0;
parameter W14TO80 = 0;
parameter W14TO81 = 0;
parameter W14TO82 = 0;
parameter W14TO83 = 0;
parameter W14TO84 = 0;
parameter W14TO85 = 0;
parameter W14TO86 = 0;
parameter W14TO87 = 0;
parameter W14TO88 = 0;
parameter W14TO89 = 0;
parameter W14TO90 = 0;
parameter W14TO91 = 0;
parameter W14TO92 = 0;
parameter W14TO93 = 0;
parameter W14TO94 = 0;
parameter W14TO95 = 0;
parameter W14TO96 = 0;
parameter W14TO97 = 0;
parameter W14TO98 = 0;
parameter W14TO99 = 0;
parameter W15TO0 = 0;
parameter W15TO1 = 0;
parameter W15TO2 = 0;
parameter W15TO3 = 0;
parameter W15TO4 = 0;
parameter W15TO5 = 0;
parameter W15TO6 = 0;
parameter W15TO7 = 0;
parameter W15TO8 = 0;
parameter W15TO9 = 0;
parameter W15TO10 = 0;
parameter W15TO11 = 0;
parameter W15TO12 = 0;
parameter W15TO13 = 0;
parameter W15TO14 = 0;
parameter W15TO15 = 0;
parameter W15TO16 = 0;
parameter W15TO17 = 0;
parameter W15TO18 = 0;
parameter W15TO19 = 0;
parameter W15TO20 = 0;
parameter W15TO21 = 0;
parameter W15TO22 = 0;
parameter W15TO23 = 0;
parameter W15TO24 = 0;
parameter W15TO25 = 0;
parameter W15TO26 = 0;
parameter W15TO27 = 0;
parameter W15TO28 = 0;
parameter W15TO29 = 0;
parameter W15TO30 = 0;
parameter W15TO31 = 0;
parameter W15TO32 = 0;
parameter W15TO33 = 0;
parameter W15TO34 = 0;
parameter W15TO35 = 0;
parameter W15TO36 = 0;
parameter W15TO37 = 0;
parameter W15TO38 = 0;
parameter W15TO39 = 0;
parameter W15TO40 = 0;
parameter W15TO41 = 0;
parameter W15TO42 = 0;
parameter W15TO43 = 0;
parameter W15TO44 = 0;
parameter W15TO45 = 0;
parameter W15TO46 = 0;
parameter W15TO47 = 0;
parameter W15TO48 = 0;
parameter W15TO49 = 0;
parameter W15TO50 = 0;
parameter W15TO51 = 0;
parameter W15TO52 = 0;
parameter W15TO53 = 0;
parameter W15TO54 = 0;
parameter W15TO55 = 0;
parameter W15TO56 = 0;
parameter W15TO57 = 0;
parameter W15TO58 = 0;
parameter W15TO59 = 0;
parameter W15TO60 = 0;
parameter W15TO61 = 0;
parameter W15TO62 = 0;
parameter W15TO63 = 0;
parameter W15TO64 = 0;
parameter W15TO65 = 0;
parameter W15TO66 = 0;
parameter W15TO67 = 0;
parameter W15TO68 = 0;
parameter W15TO69 = 0;
parameter W15TO70 = 0;
parameter W15TO71 = 0;
parameter W15TO72 = 0;
parameter W15TO73 = 0;
parameter W15TO74 = 0;
parameter W15TO75 = 0;
parameter W15TO76 = 0;
parameter W15TO77 = 0;
parameter W15TO78 = 0;
parameter W15TO79 = 0;
parameter W15TO80 = 0;
parameter W15TO81 = 0;
parameter W15TO82 = 0;
parameter W15TO83 = 0;
parameter W15TO84 = 0;
parameter W15TO85 = 0;
parameter W15TO86 = 0;
parameter W15TO87 = 0;
parameter W15TO88 = 0;
parameter W15TO89 = 0;
parameter W15TO90 = 0;
parameter W15TO91 = 0;
parameter W15TO92 = 0;
parameter W15TO93 = 0;
parameter W15TO94 = 0;
parameter W15TO95 = 0;
parameter W15TO96 = 0;
parameter W15TO97 = 0;
parameter W15TO98 = 0;
parameter W15TO99 = 0;
parameter W16TO0 = 0;
parameter W16TO1 = 0;
parameter W16TO2 = 0;
parameter W16TO3 = 0;
parameter W16TO4 = 0;
parameter W16TO5 = 0;
parameter W16TO6 = 0;
parameter W16TO7 = 0;
parameter W16TO8 = 0;
parameter W16TO9 = 0;
parameter W16TO10 = 0;
parameter W16TO11 = 0;
parameter W16TO12 = 0;
parameter W16TO13 = 0;
parameter W16TO14 = 0;
parameter W16TO15 = 0;
parameter W16TO16 = 0;
parameter W16TO17 = 0;
parameter W16TO18 = 0;
parameter W16TO19 = 0;
parameter W16TO20 = 0;
parameter W16TO21 = 0;
parameter W16TO22 = 0;
parameter W16TO23 = 0;
parameter W16TO24 = 0;
parameter W16TO25 = 0;
parameter W16TO26 = 0;
parameter W16TO27 = 0;
parameter W16TO28 = 0;
parameter W16TO29 = 0;
parameter W16TO30 = 0;
parameter W16TO31 = 0;
parameter W16TO32 = 0;
parameter W16TO33 = 0;
parameter W16TO34 = 0;
parameter W16TO35 = 0;
parameter W16TO36 = 0;
parameter W16TO37 = 0;
parameter W16TO38 = 0;
parameter W16TO39 = 0;
parameter W16TO40 = 0;
parameter W16TO41 = 0;
parameter W16TO42 = 0;
parameter W16TO43 = 0;
parameter W16TO44 = 0;
parameter W16TO45 = 0;
parameter W16TO46 = 0;
parameter W16TO47 = 0;
parameter W16TO48 = 0;
parameter W16TO49 = 0;
parameter W16TO50 = 0;
parameter W16TO51 = 0;
parameter W16TO52 = 0;
parameter W16TO53 = 0;
parameter W16TO54 = 0;
parameter W16TO55 = 0;
parameter W16TO56 = 0;
parameter W16TO57 = 0;
parameter W16TO58 = 0;
parameter W16TO59 = 0;
parameter W16TO60 = 0;
parameter W16TO61 = 0;
parameter W16TO62 = 0;
parameter W16TO63 = 0;
parameter W16TO64 = 0;
parameter W16TO65 = 0;
parameter W16TO66 = 0;
parameter W16TO67 = 0;
parameter W16TO68 = 0;
parameter W16TO69 = 0;
parameter W16TO70 = 0;
parameter W16TO71 = 0;
parameter W16TO72 = 0;
parameter W16TO73 = 0;
parameter W16TO74 = 0;
parameter W16TO75 = 0;
parameter W16TO76 = 0;
parameter W16TO77 = 0;
parameter W16TO78 = 0;
parameter W16TO79 = 0;
parameter W16TO80 = 0;
parameter W16TO81 = 0;
parameter W16TO82 = 0;
parameter W16TO83 = 0;
parameter W16TO84 = 0;
parameter W16TO85 = 0;
parameter W16TO86 = 0;
parameter W16TO87 = 0;
parameter W16TO88 = 0;
parameter W16TO89 = 0;
parameter W16TO90 = 0;
parameter W16TO91 = 0;
parameter W16TO92 = 0;
parameter W16TO93 = 0;
parameter W16TO94 = 0;
parameter W16TO95 = 0;
parameter W16TO96 = 0;
parameter W16TO97 = 0;
parameter W16TO98 = 0;
parameter W16TO99 = 0;
parameter W17TO0 = 0;
parameter W17TO1 = 0;
parameter W17TO2 = 0;
parameter W17TO3 = 0;
parameter W17TO4 = 0;
parameter W17TO5 = 0;
parameter W17TO6 = 0;
parameter W17TO7 = 0;
parameter W17TO8 = 0;
parameter W17TO9 = 0;
parameter W17TO10 = 0;
parameter W17TO11 = 0;
parameter W17TO12 = 0;
parameter W17TO13 = 0;
parameter W17TO14 = 0;
parameter W17TO15 = 0;
parameter W17TO16 = 0;
parameter W17TO17 = 0;
parameter W17TO18 = 0;
parameter W17TO19 = 0;
parameter W17TO20 = 0;
parameter W17TO21 = 0;
parameter W17TO22 = 0;
parameter W17TO23 = 0;
parameter W17TO24 = 0;
parameter W17TO25 = 0;
parameter W17TO26 = 0;
parameter W17TO27 = 0;
parameter W17TO28 = 0;
parameter W17TO29 = 0;
parameter W17TO30 = 0;
parameter W17TO31 = 0;
parameter W17TO32 = 0;
parameter W17TO33 = 0;
parameter W17TO34 = 0;
parameter W17TO35 = 0;
parameter W17TO36 = 0;
parameter W17TO37 = 0;
parameter W17TO38 = 0;
parameter W17TO39 = 0;
parameter W17TO40 = 0;
parameter W17TO41 = 0;
parameter W17TO42 = 0;
parameter W17TO43 = 0;
parameter W17TO44 = 0;
parameter W17TO45 = 0;
parameter W17TO46 = 0;
parameter W17TO47 = 0;
parameter W17TO48 = 0;
parameter W17TO49 = 0;
parameter W17TO50 = 0;
parameter W17TO51 = 0;
parameter W17TO52 = 0;
parameter W17TO53 = 0;
parameter W17TO54 = 0;
parameter W17TO55 = 0;
parameter W17TO56 = 0;
parameter W17TO57 = 0;
parameter W17TO58 = 0;
parameter W17TO59 = 0;
parameter W17TO60 = 0;
parameter W17TO61 = 0;
parameter W17TO62 = 0;
parameter W17TO63 = 0;
parameter W17TO64 = 0;
parameter W17TO65 = 0;
parameter W17TO66 = 0;
parameter W17TO67 = 0;
parameter W17TO68 = 0;
parameter W17TO69 = 0;
parameter W17TO70 = 0;
parameter W17TO71 = 0;
parameter W17TO72 = 0;
parameter W17TO73 = 0;
parameter W17TO74 = 0;
parameter W17TO75 = 0;
parameter W17TO76 = 0;
parameter W17TO77 = 0;
parameter W17TO78 = 0;
parameter W17TO79 = 0;
parameter W17TO80 = 0;
parameter W17TO81 = 0;
parameter W17TO82 = 0;
parameter W17TO83 = 0;
parameter W17TO84 = 0;
parameter W17TO85 = 0;
parameter W17TO86 = 0;
parameter W17TO87 = 0;
parameter W17TO88 = 0;
parameter W17TO89 = 0;
parameter W17TO90 = 0;
parameter W17TO91 = 0;
parameter W17TO92 = 0;
parameter W17TO93 = 0;
parameter W17TO94 = 0;
parameter W17TO95 = 0;
parameter W17TO96 = 0;
parameter W17TO97 = 0;
parameter W17TO98 = 0;
parameter W17TO99 = 0;
parameter W18TO0 = 0;
parameter W18TO1 = 0;
parameter W18TO2 = 0;
parameter W18TO3 = 0;
parameter W18TO4 = 0;
parameter W18TO5 = 0;
parameter W18TO6 = 0;
parameter W18TO7 = 0;
parameter W18TO8 = 0;
parameter W18TO9 = 0;
parameter W18TO10 = 0;
parameter W18TO11 = 0;
parameter W18TO12 = 0;
parameter W18TO13 = 0;
parameter W18TO14 = 0;
parameter W18TO15 = 0;
parameter W18TO16 = 0;
parameter W18TO17 = 0;
parameter W18TO18 = 0;
parameter W18TO19 = 0;
parameter W18TO20 = 0;
parameter W18TO21 = 0;
parameter W18TO22 = 0;
parameter W18TO23 = 0;
parameter W18TO24 = 0;
parameter W18TO25 = 0;
parameter W18TO26 = 0;
parameter W18TO27 = 0;
parameter W18TO28 = 0;
parameter W18TO29 = 0;
parameter W18TO30 = 0;
parameter W18TO31 = 0;
parameter W18TO32 = 0;
parameter W18TO33 = 0;
parameter W18TO34 = 0;
parameter W18TO35 = 0;
parameter W18TO36 = 0;
parameter W18TO37 = 0;
parameter W18TO38 = 0;
parameter W18TO39 = 0;
parameter W18TO40 = 0;
parameter W18TO41 = 0;
parameter W18TO42 = 0;
parameter W18TO43 = 0;
parameter W18TO44 = 0;
parameter W18TO45 = 0;
parameter W18TO46 = 0;
parameter W18TO47 = 0;
parameter W18TO48 = 0;
parameter W18TO49 = 0;
parameter W18TO50 = 0;
parameter W18TO51 = 0;
parameter W18TO52 = 0;
parameter W18TO53 = 0;
parameter W18TO54 = 0;
parameter W18TO55 = 0;
parameter W18TO56 = 0;
parameter W18TO57 = 0;
parameter W18TO58 = 0;
parameter W18TO59 = 0;
parameter W18TO60 = 0;
parameter W18TO61 = 0;
parameter W18TO62 = 0;
parameter W18TO63 = 0;
parameter W18TO64 = 0;
parameter W18TO65 = 0;
parameter W18TO66 = 0;
parameter W18TO67 = 0;
parameter W18TO68 = 0;
parameter W18TO69 = 0;
parameter W18TO70 = 0;
parameter W18TO71 = 0;
parameter W18TO72 = 0;
parameter W18TO73 = 0;
parameter W18TO74 = 0;
parameter W18TO75 = 0;
parameter W18TO76 = 0;
parameter W18TO77 = 0;
parameter W18TO78 = 0;
parameter W18TO79 = 0;
parameter W18TO80 = 0;
parameter W18TO81 = 0;
parameter W18TO82 = 0;
parameter W18TO83 = 0;
parameter W18TO84 = 0;
parameter W18TO85 = 0;
parameter W18TO86 = 0;
parameter W18TO87 = 0;
parameter W18TO88 = 0;
parameter W18TO89 = 0;
parameter W18TO90 = 0;
parameter W18TO91 = 0;
parameter W18TO92 = 0;
parameter W18TO93 = 0;
parameter W18TO94 = 0;
parameter W18TO95 = 0;
parameter W18TO96 = 0;
parameter W18TO97 = 0;
parameter W18TO98 = 0;
parameter W18TO99 = 0;
parameter W19TO0 = 0;
parameter W19TO1 = 0;
parameter W19TO2 = 0;
parameter W19TO3 = 0;
parameter W19TO4 = 0;
parameter W19TO5 = 0;
parameter W19TO6 = 0;
parameter W19TO7 = 0;
parameter W19TO8 = 0;
parameter W19TO9 = 0;
parameter W19TO10 = 0;
parameter W19TO11 = 0;
parameter W19TO12 = 0;
parameter W19TO13 = 0;
parameter W19TO14 = 0;
parameter W19TO15 = 0;
parameter W19TO16 = 0;
parameter W19TO17 = 0;
parameter W19TO18 = 0;
parameter W19TO19 = 0;
parameter W19TO20 = 0;
parameter W19TO21 = 0;
parameter W19TO22 = 0;
parameter W19TO23 = 0;
parameter W19TO24 = 0;
parameter W19TO25 = 0;
parameter W19TO26 = 0;
parameter W19TO27 = 0;
parameter W19TO28 = 0;
parameter W19TO29 = 0;
parameter W19TO30 = 0;
parameter W19TO31 = 0;
parameter W19TO32 = 0;
parameter W19TO33 = 0;
parameter W19TO34 = 0;
parameter W19TO35 = 0;
parameter W19TO36 = 0;
parameter W19TO37 = 0;
parameter W19TO38 = 0;
parameter W19TO39 = 0;
parameter W19TO40 = 0;
parameter W19TO41 = 0;
parameter W19TO42 = 0;
parameter W19TO43 = 0;
parameter W19TO44 = 0;
parameter W19TO45 = 0;
parameter W19TO46 = 0;
parameter W19TO47 = 0;
parameter W19TO48 = 0;
parameter W19TO49 = 0;
parameter W19TO50 = 0;
parameter W19TO51 = 0;
parameter W19TO52 = 0;
parameter W19TO53 = 0;
parameter W19TO54 = 0;
parameter W19TO55 = 0;
parameter W19TO56 = 0;
parameter W19TO57 = 0;
parameter W19TO58 = 0;
parameter W19TO59 = 0;
parameter W19TO60 = 0;
parameter W19TO61 = 0;
parameter W19TO62 = 0;
parameter W19TO63 = 0;
parameter W19TO64 = 0;
parameter W19TO65 = 0;
parameter W19TO66 = 0;
parameter W19TO67 = 0;
parameter W19TO68 = 0;
parameter W19TO69 = 0;
parameter W19TO70 = 0;
parameter W19TO71 = 0;
parameter W19TO72 = 0;
parameter W19TO73 = 0;
parameter W19TO74 = 0;
parameter W19TO75 = 0;
parameter W19TO76 = 0;
parameter W19TO77 = 0;
parameter W19TO78 = 0;
parameter W19TO79 = 0;
parameter W19TO80 = 0;
parameter W19TO81 = 0;
parameter W19TO82 = 0;
parameter W19TO83 = 0;
parameter W19TO84 = 0;
parameter W19TO85 = 0;
parameter W19TO86 = 0;
parameter W19TO87 = 0;
parameter W19TO88 = 0;
parameter W19TO89 = 0;
parameter W19TO90 = 0;
parameter W19TO91 = 0;
parameter W19TO92 = 0;
parameter W19TO93 = 0;
parameter W19TO94 = 0;
parameter W19TO95 = 0;
parameter W19TO96 = 0;
parameter W19TO97 = 0;
parameter W19TO98 = 0;
parameter W19TO99 = 0;
parameter W20TO0 = 0;
parameter W20TO1 = 0;
parameter W20TO2 = 0;
parameter W20TO3 = 0;
parameter W20TO4 = 0;
parameter W20TO5 = 0;
parameter W20TO6 = 0;
parameter W20TO7 = 0;
parameter W20TO8 = 0;
parameter W20TO9 = 0;
parameter W20TO10 = 0;
parameter W20TO11 = 0;
parameter W20TO12 = 0;
parameter W20TO13 = 0;
parameter W20TO14 = 0;
parameter W20TO15 = 0;
parameter W20TO16 = 0;
parameter W20TO17 = 0;
parameter W20TO18 = 0;
parameter W20TO19 = 0;
parameter W20TO20 = 0;
parameter W20TO21 = 0;
parameter W20TO22 = 0;
parameter W20TO23 = 0;
parameter W20TO24 = 0;
parameter W20TO25 = 0;
parameter W20TO26 = 0;
parameter W20TO27 = 0;
parameter W20TO28 = 0;
parameter W20TO29 = 0;
parameter W20TO30 = 0;
parameter W20TO31 = 0;
parameter W20TO32 = 0;
parameter W20TO33 = 0;
parameter W20TO34 = 0;
parameter W20TO35 = 0;
parameter W20TO36 = 0;
parameter W20TO37 = 0;
parameter W20TO38 = 0;
parameter W20TO39 = 0;
parameter W20TO40 = 0;
parameter W20TO41 = 0;
parameter W20TO42 = 0;
parameter W20TO43 = 0;
parameter W20TO44 = 0;
parameter W20TO45 = 0;
parameter W20TO46 = 0;
parameter W20TO47 = 0;
parameter W20TO48 = 0;
parameter W20TO49 = 0;
parameter W20TO50 = 0;
parameter W20TO51 = 0;
parameter W20TO52 = 0;
parameter W20TO53 = 0;
parameter W20TO54 = 0;
parameter W20TO55 = 0;
parameter W20TO56 = 0;
parameter W20TO57 = 0;
parameter W20TO58 = 0;
parameter W20TO59 = 0;
parameter W20TO60 = 0;
parameter W20TO61 = 0;
parameter W20TO62 = 0;
parameter W20TO63 = 0;
parameter W20TO64 = 0;
parameter W20TO65 = 0;
parameter W20TO66 = 0;
parameter W20TO67 = 0;
parameter W20TO68 = 0;
parameter W20TO69 = 0;
parameter W20TO70 = 0;
parameter W20TO71 = 0;
parameter W20TO72 = 0;
parameter W20TO73 = 0;
parameter W20TO74 = 0;
parameter W20TO75 = 0;
parameter W20TO76 = 0;
parameter W20TO77 = 0;
parameter W20TO78 = 0;
parameter W20TO79 = 0;
parameter W20TO80 = 0;
parameter W20TO81 = 0;
parameter W20TO82 = 0;
parameter W20TO83 = 0;
parameter W20TO84 = 0;
parameter W20TO85 = 0;
parameter W20TO86 = 0;
parameter W20TO87 = 0;
parameter W20TO88 = 0;
parameter W20TO89 = 0;
parameter W20TO90 = 0;
parameter W20TO91 = 0;
parameter W20TO92 = 0;
parameter W20TO93 = 0;
parameter W20TO94 = 0;
parameter W20TO95 = 0;
parameter W20TO96 = 0;
parameter W20TO97 = 0;
parameter W20TO98 = 0;
parameter W20TO99 = 0;
parameter W21TO0 = 0;
parameter W21TO1 = 0;
parameter W21TO2 = 0;
parameter W21TO3 = 0;
parameter W21TO4 = 0;
parameter W21TO5 = 0;
parameter W21TO6 = 0;
parameter W21TO7 = 0;
parameter W21TO8 = 0;
parameter W21TO9 = 0;
parameter W21TO10 = 0;
parameter W21TO11 = 0;
parameter W21TO12 = 0;
parameter W21TO13 = 0;
parameter W21TO14 = 0;
parameter W21TO15 = 0;
parameter W21TO16 = 0;
parameter W21TO17 = 0;
parameter W21TO18 = 0;
parameter W21TO19 = 0;
parameter W21TO20 = 0;
parameter W21TO21 = 0;
parameter W21TO22 = 0;
parameter W21TO23 = 0;
parameter W21TO24 = 0;
parameter W21TO25 = 0;
parameter W21TO26 = 0;
parameter W21TO27 = 0;
parameter W21TO28 = 0;
parameter W21TO29 = 0;
parameter W21TO30 = 0;
parameter W21TO31 = 0;
parameter W21TO32 = 0;
parameter W21TO33 = 0;
parameter W21TO34 = 0;
parameter W21TO35 = 0;
parameter W21TO36 = 0;
parameter W21TO37 = 0;
parameter W21TO38 = 0;
parameter W21TO39 = 0;
parameter W21TO40 = 0;
parameter W21TO41 = 0;
parameter W21TO42 = 0;
parameter W21TO43 = 0;
parameter W21TO44 = 0;
parameter W21TO45 = 0;
parameter W21TO46 = 0;
parameter W21TO47 = 0;
parameter W21TO48 = 0;
parameter W21TO49 = 0;
parameter W21TO50 = 0;
parameter W21TO51 = 0;
parameter W21TO52 = 0;
parameter W21TO53 = 0;
parameter W21TO54 = 0;
parameter W21TO55 = 0;
parameter W21TO56 = 0;
parameter W21TO57 = 0;
parameter W21TO58 = 0;
parameter W21TO59 = 0;
parameter W21TO60 = 0;
parameter W21TO61 = 0;
parameter W21TO62 = 0;
parameter W21TO63 = 0;
parameter W21TO64 = 0;
parameter W21TO65 = 0;
parameter W21TO66 = 0;
parameter W21TO67 = 0;
parameter W21TO68 = 0;
parameter W21TO69 = 0;
parameter W21TO70 = 0;
parameter W21TO71 = 0;
parameter W21TO72 = 0;
parameter W21TO73 = 0;
parameter W21TO74 = 0;
parameter W21TO75 = 0;
parameter W21TO76 = 0;
parameter W21TO77 = 0;
parameter W21TO78 = 0;
parameter W21TO79 = 0;
parameter W21TO80 = 0;
parameter W21TO81 = 0;
parameter W21TO82 = 0;
parameter W21TO83 = 0;
parameter W21TO84 = 0;
parameter W21TO85 = 0;
parameter W21TO86 = 0;
parameter W21TO87 = 0;
parameter W21TO88 = 0;
parameter W21TO89 = 0;
parameter W21TO90 = 0;
parameter W21TO91 = 0;
parameter W21TO92 = 0;
parameter W21TO93 = 0;
parameter W21TO94 = 0;
parameter W21TO95 = 0;
parameter W21TO96 = 0;
parameter W21TO97 = 0;
parameter W21TO98 = 0;
parameter W21TO99 = 0;
parameter W22TO0 = 0;
parameter W22TO1 = 0;
parameter W22TO2 = 0;
parameter W22TO3 = 0;
parameter W22TO4 = 0;
parameter W22TO5 = 0;
parameter W22TO6 = 0;
parameter W22TO7 = 0;
parameter W22TO8 = 0;
parameter W22TO9 = 0;
parameter W22TO10 = 0;
parameter W22TO11 = 0;
parameter W22TO12 = 0;
parameter W22TO13 = 0;
parameter W22TO14 = 0;
parameter W22TO15 = 0;
parameter W22TO16 = 0;
parameter W22TO17 = 0;
parameter W22TO18 = 0;
parameter W22TO19 = 0;
parameter W22TO20 = 0;
parameter W22TO21 = 0;
parameter W22TO22 = 0;
parameter W22TO23 = 0;
parameter W22TO24 = 0;
parameter W22TO25 = 0;
parameter W22TO26 = 0;
parameter W22TO27 = 0;
parameter W22TO28 = 0;
parameter W22TO29 = 0;
parameter W22TO30 = 0;
parameter W22TO31 = 0;
parameter W22TO32 = 0;
parameter W22TO33 = 0;
parameter W22TO34 = 0;
parameter W22TO35 = 0;
parameter W22TO36 = 0;
parameter W22TO37 = 0;
parameter W22TO38 = 0;
parameter W22TO39 = 0;
parameter W22TO40 = 0;
parameter W22TO41 = 0;
parameter W22TO42 = 0;
parameter W22TO43 = 0;
parameter W22TO44 = 0;
parameter W22TO45 = 0;
parameter W22TO46 = 0;
parameter W22TO47 = 0;
parameter W22TO48 = 0;
parameter W22TO49 = 0;
parameter W22TO50 = 0;
parameter W22TO51 = 0;
parameter W22TO52 = 0;
parameter W22TO53 = 0;
parameter W22TO54 = 0;
parameter W22TO55 = 0;
parameter W22TO56 = 0;
parameter W22TO57 = 0;
parameter W22TO58 = 0;
parameter W22TO59 = 0;
parameter W22TO60 = 0;
parameter W22TO61 = 0;
parameter W22TO62 = 0;
parameter W22TO63 = 0;
parameter W22TO64 = 0;
parameter W22TO65 = 0;
parameter W22TO66 = 0;
parameter W22TO67 = 0;
parameter W22TO68 = 0;
parameter W22TO69 = 0;
parameter W22TO70 = 0;
parameter W22TO71 = 0;
parameter W22TO72 = 0;
parameter W22TO73 = 0;
parameter W22TO74 = 0;
parameter W22TO75 = 0;
parameter W22TO76 = 0;
parameter W22TO77 = 0;
parameter W22TO78 = 0;
parameter W22TO79 = 0;
parameter W22TO80 = 0;
parameter W22TO81 = 0;
parameter W22TO82 = 0;
parameter W22TO83 = 0;
parameter W22TO84 = 0;
parameter W22TO85 = 0;
parameter W22TO86 = 0;
parameter W22TO87 = 0;
parameter W22TO88 = 0;
parameter W22TO89 = 0;
parameter W22TO90 = 0;
parameter W22TO91 = 0;
parameter W22TO92 = 0;
parameter W22TO93 = 0;
parameter W22TO94 = 0;
parameter W22TO95 = 0;
parameter W22TO96 = 0;
parameter W22TO97 = 0;
parameter W22TO98 = 0;
parameter W22TO99 = 0;
parameter W23TO0 = 0;
parameter W23TO1 = 0;
parameter W23TO2 = 0;
parameter W23TO3 = 0;
parameter W23TO4 = 0;
parameter W23TO5 = 0;
parameter W23TO6 = 0;
parameter W23TO7 = 0;
parameter W23TO8 = 0;
parameter W23TO9 = 0;
parameter W23TO10 = 0;
parameter W23TO11 = 0;
parameter W23TO12 = 0;
parameter W23TO13 = 0;
parameter W23TO14 = 0;
parameter W23TO15 = 0;
parameter W23TO16 = 0;
parameter W23TO17 = 0;
parameter W23TO18 = 0;
parameter W23TO19 = 0;
parameter W23TO20 = 0;
parameter W23TO21 = 0;
parameter W23TO22 = 0;
parameter W23TO23 = 0;
parameter W23TO24 = 0;
parameter W23TO25 = 0;
parameter W23TO26 = 0;
parameter W23TO27 = 0;
parameter W23TO28 = 0;
parameter W23TO29 = 0;
parameter W23TO30 = 0;
parameter W23TO31 = 0;
parameter W23TO32 = 0;
parameter W23TO33 = 0;
parameter W23TO34 = 0;
parameter W23TO35 = 0;
parameter W23TO36 = 0;
parameter W23TO37 = 0;
parameter W23TO38 = 0;
parameter W23TO39 = 0;
parameter W23TO40 = 0;
parameter W23TO41 = 0;
parameter W23TO42 = 0;
parameter W23TO43 = 0;
parameter W23TO44 = 0;
parameter W23TO45 = 0;
parameter W23TO46 = 0;
parameter W23TO47 = 0;
parameter W23TO48 = 0;
parameter W23TO49 = 0;
parameter W23TO50 = 0;
parameter W23TO51 = 0;
parameter W23TO52 = 0;
parameter W23TO53 = 0;
parameter W23TO54 = 0;
parameter W23TO55 = 0;
parameter W23TO56 = 0;
parameter W23TO57 = 0;
parameter W23TO58 = 0;
parameter W23TO59 = 0;
parameter W23TO60 = 0;
parameter W23TO61 = 0;
parameter W23TO62 = 0;
parameter W23TO63 = 0;
parameter W23TO64 = 0;
parameter W23TO65 = 0;
parameter W23TO66 = 0;
parameter W23TO67 = 0;
parameter W23TO68 = 0;
parameter W23TO69 = 0;
parameter W23TO70 = 0;
parameter W23TO71 = 0;
parameter W23TO72 = 0;
parameter W23TO73 = 0;
parameter W23TO74 = 0;
parameter W23TO75 = 0;
parameter W23TO76 = 0;
parameter W23TO77 = 0;
parameter W23TO78 = 0;
parameter W23TO79 = 0;
parameter W23TO80 = 0;
parameter W23TO81 = 0;
parameter W23TO82 = 0;
parameter W23TO83 = 0;
parameter W23TO84 = 0;
parameter W23TO85 = 0;
parameter W23TO86 = 0;
parameter W23TO87 = 0;
parameter W23TO88 = 0;
parameter W23TO89 = 0;
parameter W23TO90 = 0;
parameter W23TO91 = 0;
parameter W23TO92 = 0;
parameter W23TO93 = 0;
parameter W23TO94 = 0;
parameter W23TO95 = 0;
parameter W23TO96 = 0;
parameter W23TO97 = 0;
parameter W23TO98 = 0;
parameter W23TO99 = 0;
parameter W24TO0 = 0;
parameter W24TO1 = 0;
parameter W24TO2 = 0;
parameter W24TO3 = 0;
parameter W24TO4 = 0;
parameter W24TO5 = 0;
parameter W24TO6 = 0;
parameter W24TO7 = 0;
parameter W24TO8 = 0;
parameter W24TO9 = 0;
parameter W24TO10 = 0;
parameter W24TO11 = 0;
parameter W24TO12 = 0;
parameter W24TO13 = 0;
parameter W24TO14 = 0;
parameter W24TO15 = 0;
parameter W24TO16 = 0;
parameter W24TO17 = 0;
parameter W24TO18 = 0;
parameter W24TO19 = 0;
parameter W24TO20 = 0;
parameter W24TO21 = 0;
parameter W24TO22 = 0;
parameter W24TO23 = 0;
parameter W24TO24 = 0;
parameter W24TO25 = 0;
parameter W24TO26 = 0;
parameter W24TO27 = 0;
parameter W24TO28 = 0;
parameter W24TO29 = 0;
parameter W24TO30 = 0;
parameter W24TO31 = 0;
parameter W24TO32 = 0;
parameter W24TO33 = 0;
parameter W24TO34 = 0;
parameter W24TO35 = 0;
parameter W24TO36 = 0;
parameter W24TO37 = 0;
parameter W24TO38 = 0;
parameter W24TO39 = 0;
parameter W24TO40 = 0;
parameter W24TO41 = 0;
parameter W24TO42 = 0;
parameter W24TO43 = 0;
parameter W24TO44 = 0;
parameter W24TO45 = 0;
parameter W24TO46 = 0;
parameter W24TO47 = 0;
parameter W24TO48 = 0;
parameter W24TO49 = 0;
parameter W24TO50 = 0;
parameter W24TO51 = 0;
parameter W24TO52 = 0;
parameter W24TO53 = 0;
parameter W24TO54 = 0;
parameter W24TO55 = 0;
parameter W24TO56 = 0;
parameter W24TO57 = 0;
parameter W24TO58 = 0;
parameter W24TO59 = 0;
parameter W24TO60 = 0;
parameter W24TO61 = 0;
parameter W24TO62 = 0;
parameter W24TO63 = 0;
parameter W24TO64 = 0;
parameter W24TO65 = 0;
parameter W24TO66 = 0;
parameter W24TO67 = 0;
parameter W24TO68 = 0;
parameter W24TO69 = 0;
parameter W24TO70 = 0;
parameter W24TO71 = 0;
parameter W24TO72 = 0;
parameter W24TO73 = 0;
parameter W24TO74 = 0;
parameter W24TO75 = 0;
parameter W24TO76 = 0;
parameter W24TO77 = 0;
parameter W24TO78 = 0;
parameter W24TO79 = 0;
parameter W24TO80 = 0;
parameter W24TO81 = 0;
parameter W24TO82 = 0;
parameter W24TO83 = 0;
parameter W24TO84 = 0;
parameter W24TO85 = 0;
parameter W24TO86 = 0;
parameter W24TO87 = 0;
parameter W24TO88 = 0;
parameter W24TO89 = 0;
parameter W24TO90 = 0;
parameter W24TO91 = 0;
parameter W24TO92 = 0;
parameter W24TO93 = 0;
parameter W24TO94 = 0;
parameter W24TO95 = 0;
parameter W24TO96 = 0;
parameter W24TO97 = 0;
parameter W24TO98 = 0;
parameter W24TO99 = 0;
parameter W25TO0 = 0;
parameter W25TO1 = 0;
parameter W25TO2 = 0;
parameter W25TO3 = 0;
parameter W25TO4 = 0;
parameter W25TO5 = 0;
parameter W25TO6 = 0;
parameter W25TO7 = 0;
parameter W25TO8 = 0;
parameter W25TO9 = 0;
parameter W25TO10 = 0;
parameter W25TO11 = 0;
parameter W25TO12 = 0;
parameter W25TO13 = 0;
parameter W25TO14 = 0;
parameter W25TO15 = 0;
parameter W25TO16 = 0;
parameter W25TO17 = 0;
parameter W25TO18 = 0;
parameter W25TO19 = 0;
parameter W25TO20 = 0;
parameter W25TO21 = 0;
parameter W25TO22 = 0;
parameter W25TO23 = 0;
parameter W25TO24 = 0;
parameter W25TO25 = 0;
parameter W25TO26 = 0;
parameter W25TO27 = 0;
parameter W25TO28 = 0;
parameter W25TO29 = 0;
parameter W25TO30 = 0;
parameter W25TO31 = 0;
parameter W25TO32 = 0;
parameter W25TO33 = 0;
parameter W25TO34 = 0;
parameter W25TO35 = 0;
parameter W25TO36 = 0;
parameter W25TO37 = 0;
parameter W25TO38 = 0;
parameter W25TO39 = 0;
parameter W25TO40 = 0;
parameter W25TO41 = 0;
parameter W25TO42 = 0;
parameter W25TO43 = 0;
parameter W25TO44 = 0;
parameter W25TO45 = 0;
parameter W25TO46 = 0;
parameter W25TO47 = 0;
parameter W25TO48 = 0;
parameter W25TO49 = 0;
parameter W25TO50 = 0;
parameter W25TO51 = 0;
parameter W25TO52 = 0;
parameter W25TO53 = 0;
parameter W25TO54 = 0;
parameter W25TO55 = 0;
parameter W25TO56 = 0;
parameter W25TO57 = 0;
parameter W25TO58 = 0;
parameter W25TO59 = 0;
parameter W25TO60 = 0;
parameter W25TO61 = 0;
parameter W25TO62 = 0;
parameter W25TO63 = 0;
parameter W25TO64 = 0;
parameter W25TO65 = 0;
parameter W25TO66 = 0;
parameter W25TO67 = 0;
parameter W25TO68 = 0;
parameter W25TO69 = 0;
parameter W25TO70 = 0;
parameter W25TO71 = 0;
parameter W25TO72 = 0;
parameter W25TO73 = 0;
parameter W25TO74 = 0;
parameter W25TO75 = 0;
parameter W25TO76 = 0;
parameter W25TO77 = 0;
parameter W25TO78 = 0;
parameter W25TO79 = 0;
parameter W25TO80 = 0;
parameter W25TO81 = 0;
parameter W25TO82 = 0;
parameter W25TO83 = 0;
parameter W25TO84 = 0;
parameter W25TO85 = 0;
parameter W25TO86 = 0;
parameter W25TO87 = 0;
parameter W25TO88 = 0;
parameter W25TO89 = 0;
parameter W25TO90 = 0;
parameter W25TO91 = 0;
parameter W25TO92 = 0;
parameter W25TO93 = 0;
parameter W25TO94 = 0;
parameter W25TO95 = 0;
parameter W25TO96 = 0;
parameter W25TO97 = 0;
parameter W25TO98 = 0;
parameter W25TO99 = 0;
parameter W26TO0 = 0;
parameter W26TO1 = 0;
parameter W26TO2 = 0;
parameter W26TO3 = 0;
parameter W26TO4 = 0;
parameter W26TO5 = 0;
parameter W26TO6 = 0;
parameter W26TO7 = 0;
parameter W26TO8 = 0;
parameter W26TO9 = 0;
parameter W26TO10 = 0;
parameter W26TO11 = 0;
parameter W26TO12 = 0;
parameter W26TO13 = 0;
parameter W26TO14 = 0;
parameter W26TO15 = 0;
parameter W26TO16 = 0;
parameter W26TO17 = 0;
parameter W26TO18 = 0;
parameter W26TO19 = 0;
parameter W26TO20 = 0;
parameter W26TO21 = 0;
parameter W26TO22 = 0;
parameter W26TO23 = 0;
parameter W26TO24 = 0;
parameter W26TO25 = 0;
parameter W26TO26 = 0;
parameter W26TO27 = 0;
parameter W26TO28 = 0;
parameter W26TO29 = 0;
parameter W26TO30 = 0;
parameter W26TO31 = 0;
parameter W26TO32 = 0;
parameter W26TO33 = 0;
parameter W26TO34 = 0;
parameter W26TO35 = 0;
parameter W26TO36 = 0;
parameter W26TO37 = 0;
parameter W26TO38 = 0;
parameter W26TO39 = 0;
parameter W26TO40 = 0;
parameter W26TO41 = 0;
parameter W26TO42 = 0;
parameter W26TO43 = 0;
parameter W26TO44 = 0;
parameter W26TO45 = 0;
parameter W26TO46 = 0;
parameter W26TO47 = 0;
parameter W26TO48 = 0;
parameter W26TO49 = 0;
parameter W26TO50 = 0;
parameter W26TO51 = 0;
parameter W26TO52 = 0;
parameter W26TO53 = 0;
parameter W26TO54 = 0;
parameter W26TO55 = 0;
parameter W26TO56 = 0;
parameter W26TO57 = 0;
parameter W26TO58 = 0;
parameter W26TO59 = 0;
parameter W26TO60 = 0;
parameter W26TO61 = 0;
parameter W26TO62 = 0;
parameter W26TO63 = 0;
parameter W26TO64 = 0;
parameter W26TO65 = 0;
parameter W26TO66 = 0;
parameter W26TO67 = 0;
parameter W26TO68 = 0;
parameter W26TO69 = 0;
parameter W26TO70 = 0;
parameter W26TO71 = 0;
parameter W26TO72 = 0;
parameter W26TO73 = 0;
parameter W26TO74 = 0;
parameter W26TO75 = 0;
parameter W26TO76 = 0;
parameter W26TO77 = 0;
parameter W26TO78 = 0;
parameter W26TO79 = 0;
parameter W26TO80 = 0;
parameter W26TO81 = 0;
parameter W26TO82 = 0;
parameter W26TO83 = 0;
parameter W26TO84 = 0;
parameter W26TO85 = 0;
parameter W26TO86 = 0;
parameter W26TO87 = 0;
parameter W26TO88 = 0;
parameter W26TO89 = 0;
parameter W26TO90 = 0;
parameter W26TO91 = 0;
parameter W26TO92 = 0;
parameter W26TO93 = 0;
parameter W26TO94 = 0;
parameter W26TO95 = 0;
parameter W26TO96 = 0;
parameter W26TO97 = 0;
parameter W26TO98 = 0;
parameter W26TO99 = 0;
parameter W27TO0 = 0;
parameter W27TO1 = 0;
parameter W27TO2 = 0;
parameter W27TO3 = 0;
parameter W27TO4 = 0;
parameter W27TO5 = 0;
parameter W27TO6 = 0;
parameter W27TO7 = 0;
parameter W27TO8 = 0;
parameter W27TO9 = 0;
parameter W27TO10 = 0;
parameter W27TO11 = 0;
parameter W27TO12 = 0;
parameter W27TO13 = 0;
parameter W27TO14 = 0;
parameter W27TO15 = 0;
parameter W27TO16 = 0;
parameter W27TO17 = 0;
parameter W27TO18 = 0;
parameter W27TO19 = 0;
parameter W27TO20 = 0;
parameter W27TO21 = 0;
parameter W27TO22 = 0;
parameter W27TO23 = 0;
parameter W27TO24 = 0;
parameter W27TO25 = 0;
parameter W27TO26 = 0;
parameter W27TO27 = 0;
parameter W27TO28 = 0;
parameter W27TO29 = 0;
parameter W27TO30 = 0;
parameter W27TO31 = 0;
parameter W27TO32 = 0;
parameter W27TO33 = 0;
parameter W27TO34 = 0;
parameter W27TO35 = 0;
parameter W27TO36 = 0;
parameter W27TO37 = 0;
parameter W27TO38 = 0;
parameter W27TO39 = 0;
parameter W27TO40 = 0;
parameter W27TO41 = 0;
parameter W27TO42 = 0;
parameter W27TO43 = 0;
parameter W27TO44 = 0;
parameter W27TO45 = 0;
parameter W27TO46 = 0;
parameter W27TO47 = 0;
parameter W27TO48 = 0;
parameter W27TO49 = 0;
parameter W27TO50 = 0;
parameter W27TO51 = 0;
parameter W27TO52 = 0;
parameter W27TO53 = 0;
parameter W27TO54 = 0;
parameter W27TO55 = 0;
parameter W27TO56 = 0;
parameter W27TO57 = 0;
parameter W27TO58 = 0;
parameter W27TO59 = 0;
parameter W27TO60 = 0;
parameter W27TO61 = 0;
parameter W27TO62 = 0;
parameter W27TO63 = 0;
parameter W27TO64 = 0;
parameter W27TO65 = 0;
parameter W27TO66 = 0;
parameter W27TO67 = 0;
parameter W27TO68 = 0;
parameter W27TO69 = 0;
parameter W27TO70 = 0;
parameter W27TO71 = 0;
parameter W27TO72 = 0;
parameter W27TO73 = 0;
parameter W27TO74 = 0;
parameter W27TO75 = 0;
parameter W27TO76 = 0;
parameter W27TO77 = 0;
parameter W27TO78 = 0;
parameter W27TO79 = 0;
parameter W27TO80 = 0;
parameter W27TO81 = 0;
parameter W27TO82 = 0;
parameter W27TO83 = 0;
parameter W27TO84 = 0;
parameter W27TO85 = 0;
parameter W27TO86 = 0;
parameter W27TO87 = 0;
parameter W27TO88 = 0;
parameter W27TO89 = 0;
parameter W27TO90 = 0;
parameter W27TO91 = 0;
parameter W27TO92 = 0;
parameter W27TO93 = 0;
parameter W27TO94 = 0;
parameter W27TO95 = 0;
parameter W27TO96 = 0;
parameter W27TO97 = 0;
parameter W27TO98 = 0;
parameter W27TO99 = 0;
parameter W28TO0 = 0;
parameter W28TO1 = 0;
parameter W28TO2 = 0;
parameter W28TO3 = 0;
parameter W28TO4 = 0;
parameter W28TO5 = 0;
parameter W28TO6 = 0;
parameter W28TO7 = 0;
parameter W28TO8 = 0;
parameter W28TO9 = 0;
parameter W28TO10 = 0;
parameter W28TO11 = 0;
parameter W28TO12 = 0;
parameter W28TO13 = 0;
parameter W28TO14 = 0;
parameter W28TO15 = 0;
parameter W28TO16 = 0;
parameter W28TO17 = 0;
parameter W28TO18 = 0;
parameter W28TO19 = 0;
parameter W28TO20 = 0;
parameter W28TO21 = 0;
parameter W28TO22 = 0;
parameter W28TO23 = 0;
parameter W28TO24 = 0;
parameter W28TO25 = 0;
parameter W28TO26 = 0;
parameter W28TO27 = 0;
parameter W28TO28 = 0;
parameter W28TO29 = 0;
parameter W28TO30 = 0;
parameter W28TO31 = 0;
parameter W28TO32 = 0;
parameter W28TO33 = 0;
parameter W28TO34 = 0;
parameter W28TO35 = 0;
parameter W28TO36 = 0;
parameter W28TO37 = 0;
parameter W28TO38 = 0;
parameter W28TO39 = 0;
parameter W28TO40 = 0;
parameter W28TO41 = 0;
parameter W28TO42 = 0;
parameter W28TO43 = 0;
parameter W28TO44 = 0;
parameter W28TO45 = 0;
parameter W28TO46 = 0;
parameter W28TO47 = 0;
parameter W28TO48 = 0;
parameter W28TO49 = 0;
parameter W28TO50 = 0;
parameter W28TO51 = 0;
parameter W28TO52 = 0;
parameter W28TO53 = 0;
parameter W28TO54 = 0;
parameter W28TO55 = 0;
parameter W28TO56 = 0;
parameter W28TO57 = 0;
parameter W28TO58 = 0;
parameter W28TO59 = 0;
parameter W28TO60 = 0;
parameter W28TO61 = 0;
parameter W28TO62 = 0;
parameter W28TO63 = 0;
parameter W28TO64 = 0;
parameter W28TO65 = 0;
parameter W28TO66 = 0;
parameter W28TO67 = 0;
parameter W28TO68 = 0;
parameter W28TO69 = 0;
parameter W28TO70 = 0;
parameter W28TO71 = 0;
parameter W28TO72 = 0;
parameter W28TO73 = 0;
parameter W28TO74 = 0;
parameter W28TO75 = 0;
parameter W28TO76 = 0;
parameter W28TO77 = 0;
parameter W28TO78 = 0;
parameter W28TO79 = 0;
parameter W28TO80 = 0;
parameter W28TO81 = 0;
parameter W28TO82 = 0;
parameter W28TO83 = 0;
parameter W28TO84 = 0;
parameter W28TO85 = 0;
parameter W28TO86 = 0;
parameter W28TO87 = 0;
parameter W28TO88 = 0;
parameter W28TO89 = 0;
parameter W28TO90 = 0;
parameter W28TO91 = 0;
parameter W28TO92 = 0;
parameter W28TO93 = 0;
parameter W28TO94 = 0;
parameter W28TO95 = 0;
parameter W28TO96 = 0;
parameter W28TO97 = 0;
parameter W28TO98 = 0;
parameter W28TO99 = 0;
parameter W29TO0 = 0;
parameter W29TO1 = 0;
parameter W29TO2 = 0;
parameter W29TO3 = 0;
parameter W29TO4 = 0;
parameter W29TO5 = 0;
parameter W29TO6 = 0;
parameter W29TO7 = 0;
parameter W29TO8 = 0;
parameter W29TO9 = 0;
parameter W29TO10 = 0;
parameter W29TO11 = 0;
parameter W29TO12 = 0;
parameter W29TO13 = 0;
parameter W29TO14 = 0;
parameter W29TO15 = 0;
parameter W29TO16 = 0;
parameter W29TO17 = 0;
parameter W29TO18 = 0;
parameter W29TO19 = 0;
parameter W29TO20 = 0;
parameter W29TO21 = 0;
parameter W29TO22 = 0;
parameter W29TO23 = 0;
parameter W29TO24 = 0;
parameter W29TO25 = 0;
parameter W29TO26 = 0;
parameter W29TO27 = 0;
parameter W29TO28 = 0;
parameter W29TO29 = 0;
parameter W29TO30 = 0;
parameter W29TO31 = 0;
parameter W29TO32 = 0;
parameter W29TO33 = 0;
parameter W29TO34 = 0;
parameter W29TO35 = 0;
parameter W29TO36 = 0;
parameter W29TO37 = 0;
parameter W29TO38 = 0;
parameter W29TO39 = 0;
parameter W29TO40 = 0;
parameter W29TO41 = 0;
parameter W29TO42 = 0;
parameter W29TO43 = 0;
parameter W29TO44 = 0;
parameter W29TO45 = 0;
parameter W29TO46 = 0;
parameter W29TO47 = 0;
parameter W29TO48 = 0;
parameter W29TO49 = 0;
parameter W29TO50 = 0;
parameter W29TO51 = 0;
parameter W29TO52 = 0;
parameter W29TO53 = 0;
parameter W29TO54 = 0;
parameter W29TO55 = 0;
parameter W29TO56 = 0;
parameter W29TO57 = 0;
parameter W29TO58 = 0;
parameter W29TO59 = 0;
parameter W29TO60 = 0;
parameter W29TO61 = 0;
parameter W29TO62 = 0;
parameter W29TO63 = 0;
parameter W29TO64 = 0;
parameter W29TO65 = 0;
parameter W29TO66 = 0;
parameter W29TO67 = 0;
parameter W29TO68 = 0;
parameter W29TO69 = 0;
parameter W29TO70 = 0;
parameter W29TO71 = 0;
parameter W29TO72 = 0;
parameter W29TO73 = 0;
parameter W29TO74 = 0;
parameter W29TO75 = 0;
parameter W29TO76 = 0;
parameter W29TO77 = 0;
parameter W29TO78 = 0;
parameter W29TO79 = 0;
parameter W29TO80 = 0;
parameter W29TO81 = 0;
parameter W29TO82 = 0;
parameter W29TO83 = 0;
parameter W29TO84 = 0;
parameter W29TO85 = 0;
parameter W29TO86 = 0;
parameter W29TO87 = 0;
parameter W29TO88 = 0;
parameter W29TO89 = 0;
parameter W29TO90 = 0;
parameter W29TO91 = 0;
parameter W29TO92 = 0;
parameter W29TO93 = 0;
parameter W29TO94 = 0;
parameter W29TO95 = 0;
parameter W29TO96 = 0;
parameter W29TO97 = 0;
parameter W29TO98 = 0;
parameter W29TO99 = 0;
parameter W30TO0 = 0;
parameter W30TO1 = 0;
parameter W30TO2 = 0;
parameter W30TO3 = 0;
parameter W30TO4 = 0;
parameter W30TO5 = 0;
parameter W30TO6 = 0;
parameter W30TO7 = 0;
parameter W30TO8 = 0;
parameter W30TO9 = 0;
parameter W30TO10 = 0;
parameter W30TO11 = 0;
parameter W30TO12 = 0;
parameter W30TO13 = 0;
parameter W30TO14 = 0;
parameter W30TO15 = 0;
parameter W30TO16 = 0;
parameter W30TO17 = 0;
parameter W30TO18 = 0;
parameter W30TO19 = 0;
parameter W30TO20 = 0;
parameter W30TO21 = 0;
parameter W30TO22 = 0;
parameter W30TO23 = 0;
parameter W30TO24 = 0;
parameter W30TO25 = 0;
parameter W30TO26 = 0;
parameter W30TO27 = 0;
parameter W30TO28 = 0;
parameter W30TO29 = 0;
parameter W30TO30 = 0;
parameter W30TO31 = 0;
parameter W30TO32 = 0;
parameter W30TO33 = 0;
parameter W30TO34 = 0;
parameter W30TO35 = 0;
parameter W30TO36 = 0;
parameter W30TO37 = 0;
parameter W30TO38 = 0;
parameter W30TO39 = 0;
parameter W30TO40 = 0;
parameter W30TO41 = 0;
parameter W30TO42 = 0;
parameter W30TO43 = 0;
parameter W30TO44 = 0;
parameter W30TO45 = 0;
parameter W30TO46 = 0;
parameter W30TO47 = 0;
parameter W30TO48 = 0;
parameter W30TO49 = 0;
parameter W30TO50 = 0;
parameter W30TO51 = 0;
parameter W30TO52 = 0;
parameter W30TO53 = 0;
parameter W30TO54 = 0;
parameter W30TO55 = 0;
parameter W30TO56 = 0;
parameter W30TO57 = 0;
parameter W30TO58 = 0;
parameter W30TO59 = 0;
parameter W30TO60 = 0;
parameter W30TO61 = 0;
parameter W30TO62 = 0;
parameter W30TO63 = 0;
parameter W30TO64 = 0;
parameter W30TO65 = 0;
parameter W30TO66 = 0;
parameter W30TO67 = 0;
parameter W30TO68 = 0;
parameter W30TO69 = 0;
parameter W30TO70 = 0;
parameter W30TO71 = 0;
parameter W30TO72 = 0;
parameter W30TO73 = 0;
parameter W30TO74 = 0;
parameter W30TO75 = 0;
parameter W30TO76 = 0;
parameter W30TO77 = 0;
parameter W30TO78 = 0;
parameter W30TO79 = 0;
parameter W30TO80 = 0;
parameter W30TO81 = 0;
parameter W30TO82 = 0;
parameter W30TO83 = 0;
parameter W30TO84 = 0;
parameter W30TO85 = 0;
parameter W30TO86 = 0;
parameter W30TO87 = 0;
parameter W30TO88 = 0;
parameter W30TO89 = 0;
parameter W30TO90 = 0;
parameter W30TO91 = 0;
parameter W30TO92 = 0;
parameter W30TO93 = 0;
parameter W30TO94 = 0;
parameter W30TO95 = 0;
parameter W30TO96 = 0;
parameter W30TO97 = 0;
parameter W30TO98 = 0;
parameter W30TO99 = 0;
parameter W31TO0 = 0;
parameter W31TO1 = 0;
parameter W31TO2 = 0;
parameter W31TO3 = 0;
parameter W31TO4 = 0;
parameter W31TO5 = 0;
parameter W31TO6 = 0;
parameter W31TO7 = 0;
parameter W31TO8 = 0;
parameter W31TO9 = 0;
parameter W31TO10 = 0;
parameter W31TO11 = 0;
parameter W31TO12 = 0;
parameter W31TO13 = 0;
parameter W31TO14 = 0;
parameter W31TO15 = 0;
parameter W31TO16 = 0;
parameter W31TO17 = 0;
parameter W31TO18 = 0;
parameter W31TO19 = 0;
parameter W31TO20 = 0;
parameter W31TO21 = 0;
parameter W31TO22 = 0;
parameter W31TO23 = 0;
parameter W31TO24 = 0;
parameter W31TO25 = 0;
parameter W31TO26 = 0;
parameter W31TO27 = 0;
parameter W31TO28 = 0;
parameter W31TO29 = 0;
parameter W31TO30 = 0;
parameter W31TO31 = 0;
parameter W31TO32 = 0;
parameter W31TO33 = 0;
parameter W31TO34 = 0;
parameter W31TO35 = 0;
parameter W31TO36 = 0;
parameter W31TO37 = 0;
parameter W31TO38 = 0;
parameter W31TO39 = 0;
parameter W31TO40 = 0;
parameter W31TO41 = 0;
parameter W31TO42 = 0;
parameter W31TO43 = 0;
parameter W31TO44 = 0;
parameter W31TO45 = 0;
parameter W31TO46 = 0;
parameter W31TO47 = 0;
parameter W31TO48 = 0;
parameter W31TO49 = 0;
parameter W31TO50 = 0;
parameter W31TO51 = 0;
parameter W31TO52 = 0;
parameter W31TO53 = 0;
parameter W31TO54 = 0;
parameter W31TO55 = 0;
parameter W31TO56 = 0;
parameter W31TO57 = 0;
parameter W31TO58 = 0;
parameter W31TO59 = 0;
parameter W31TO60 = 0;
parameter W31TO61 = 0;
parameter W31TO62 = 0;
parameter W31TO63 = 0;
parameter W31TO64 = 0;
parameter W31TO65 = 0;
parameter W31TO66 = 0;
parameter W31TO67 = 0;
parameter W31TO68 = 0;
parameter W31TO69 = 0;
parameter W31TO70 = 0;
parameter W31TO71 = 0;
parameter W31TO72 = 0;
parameter W31TO73 = 0;
parameter W31TO74 = 0;
parameter W31TO75 = 0;
parameter W31TO76 = 0;
parameter W31TO77 = 0;
parameter W31TO78 = 0;
parameter W31TO79 = 0;
parameter W31TO80 = 0;
parameter W31TO81 = 0;
parameter W31TO82 = 0;
parameter W31TO83 = 0;
parameter W31TO84 = 0;
parameter W31TO85 = 0;
parameter W31TO86 = 0;
parameter W31TO87 = 0;
parameter W31TO88 = 0;
parameter W31TO89 = 0;
parameter W31TO90 = 0;
parameter W31TO91 = 0;
parameter W31TO92 = 0;
parameter W31TO93 = 0;
parameter W31TO94 = 0;
parameter W31TO95 = 0;
parameter W31TO96 = 0;
parameter W31TO97 = 0;
parameter W31TO98 = 0;
parameter W31TO99 = 0;
parameter W32TO0 = 0;
parameter W32TO1 = 0;
parameter W32TO2 = 0;
parameter W32TO3 = 0;
parameter W32TO4 = 0;
parameter W32TO5 = 0;
parameter W32TO6 = 0;
parameter W32TO7 = 0;
parameter W32TO8 = 0;
parameter W32TO9 = 0;
parameter W32TO10 = 0;
parameter W32TO11 = 0;
parameter W32TO12 = 0;
parameter W32TO13 = 0;
parameter W32TO14 = 0;
parameter W32TO15 = 0;
parameter W32TO16 = 0;
parameter W32TO17 = 0;
parameter W32TO18 = 0;
parameter W32TO19 = 0;
parameter W32TO20 = 0;
parameter W32TO21 = 0;
parameter W32TO22 = 0;
parameter W32TO23 = 0;
parameter W32TO24 = 0;
parameter W32TO25 = 0;
parameter W32TO26 = 0;
parameter W32TO27 = 0;
parameter W32TO28 = 0;
parameter W32TO29 = 0;
parameter W32TO30 = 0;
parameter W32TO31 = 0;
parameter W32TO32 = 0;
parameter W32TO33 = 0;
parameter W32TO34 = 0;
parameter W32TO35 = 0;
parameter W32TO36 = 0;
parameter W32TO37 = 0;
parameter W32TO38 = 0;
parameter W32TO39 = 0;
parameter W32TO40 = 0;
parameter W32TO41 = 0;
parameter W32TO42 = 0;
parameter W32TO43 = 0;
parameter W32TO44 = 0;
parameter W32TO45 = 0;
parameter W32TO46 = 0;
parameter W32TO47 = 0;
parameter W32TO48 = 0;
parameter W32TO49 = 0;
parameter W32TO50 = 0;
parameter W32TO51 = 0;
parameter W32TO52 = 0;
parameter W32TO53 = 0;
parameter W32TO54 = 0;
parameter W32TO55 = 0;
parameter W32TO56 = 0;
parameter W32TO57 = 0;
parameter W32TO58 = 0;
parameter W32TO59 = 0;
parameter W32TO60 = 0;
parameter W32TO61 = 0;
parameter W32TO62 = 0;
parameter W32TO63 = 0;
parameter W32TO64 = 0;
parameter W32TO65 = 0;
parameter W32TO66 = 0;
parameter W32TO67 = 0;
parameter W32TO68 = 0;
parameter W32TO69 = 0;
parameter W32TO70 = 0;
parameter W32TO71 = 0;
parameter W32TO72 = 0;
parameter W32TO73 = 0;
parameter W32TO74 = 0;
parameter W32TO75 = 0;
parameter W32TO76 = 0;
parameter W32TO77 = 0;
parameter W32TO78 = 0;
parameter W32TO79 = 0;
parameter W32TO80 = 0;
parameter W32TO81 = 0;
parameter W32TO82 = 0;
parameter W32TO83 = 0;
parameter W32TO84 = 0;
parameter W32TO85 = 0;
parameter W32TO86 = 0;
parameter W32TO87 = 0;
parameter W32TO88 = 0;
parameter W32TO89 = 0;
parameter W32TO90 = 0;
parameter W32TO91 = 0;
parameter W32TO92 = 0;
parameter W32TO93 = 0;
parameter W32TO94 = 0;
parameter W32TO95 = 0;
parameter W32TO96 = 0;
parameter W32TO97 = 0;
parameter W32TO98 = 0;
parameter W32TO99 = 0;
parameter W33TO0 = 0;
parameter W33TO1 = 0;
parameter W33TO2 = 0;
parameter W33TO3 = 0;
parameter W33TO4 = 0;
parameter W33TO5 = 0;
parameter W33TO6 = 0;
parameter W33TO7 = 0;
parameter W33TO8 = 0;
parameter W33TO9 = 0;
parameter W33TO10 = 0;
parameter W33TO11 = 0;
parameter W33TO12 = 0;
parameter W33TO13 = 0;
parameter W33TO14 = 0;
parameter W33TO15 = 0;
parameter W33TO16 = 0;
parameter W33TO17 = 0;
parameter W33TO18 = 0;
parameter W33TO19 = 0;
parameter W33TO20 = 0;
parameter W33TO21 = 0;
parameter W33TO22 = 0;
parameter W33TO23 = 0;
parameter W33TO24 = 0;
parameter W33TO25 = 0;
parameter W33TO26 = 0;
parameter W33TO27 = 0;
parameter W33TO28 = 0;
parameter W33TO29 = 0;
parameter W33TO30 = 0;
parameter W33TO31 = 0;
parameter W33TO32 = 0;
parameter W33TO33 = 0;
parameter W33TO34 = 0;
parameter W33TO35 = 0;
parameter W33TO36 = 0;
parameter W33TO37 = 0;
parameter W33TO38 = 0;
parameter W33TO39 = 0;
parameter W33TO40 = 0;
parameter W33TO41 = 0;
parameter W33TO42 = 0;
parameter W33TO43 = 0;
parameter W33TO44 = 0;
parameter W33TO45 = 0;
parameter W33TO46 = 0;
parameter W33TO47 = 0;
parameter W33TO48 = 0;
parameter W33TO49 = 0;
parameter W33TO50 = 0;
parameter W33TO51 = 0;
parameter W33TO52 = 0;
parameter W33TO53 = 0;
parameter W33TO54 = 0;
parameter W33TO55 = 0;
parameter W33TO56 = 0;
parameter W33TO57 = 0;
parameter W33TO58 = 0;
parameter W33TO59 = 0;
parameter W33TO60 = 0;
parameter W33TO61 = 0;
parameter W33TO62 = 0;
parameter W33TO63 = 0;
parameter W33TO64 = 0;
parameter W33TO65 = 0;
parameter W33TO66 = 0;
parameter W33TO67 = 0;
parameter W33TO68 = 0;
parameter W33TO69 = 0;
parameter W33TO70 = 0;
parameter W33TO71 = 0;
parameter W33TO72 = 0;
parameter W33TO73 = 0;
parameter W33TO74 = 0;
parameter W33TO75 = 0;
parameter W33TO76 = 0;
parameter W33TO77 = 0;
parameter W33TO78 = 0;
parameter W33TO79 = 0;
parameter W33TO80 = 0;
parameter W33TO81 = 0;
parameter W33TO82 = 0;
parameter W33TO83 = 0;
parameter W33TO84 = 0;
parameter W33TO85 = 0;
parameter W33TO86 = 0;
parameter W33TO87 = 0;
parameter W33TO88 = 0;
parameter W33TO89 = 0;
parameter W33TO90 = 0;
parameter W33TO91 = 0;
parameter W33TO92 = 0;
parameter W33TO93 = 0;
parameter W33TO94 = 0;
parameter W33TO95 = 0;
parameter W33TO96 = 0;
parameter W33TO97 = 0;
parameter W33TO98 = 0;
parameter W33TO99 = 0;
parameter W34TO0 = 0;
parameter W34TO1 = 0;
parameter W34TO2 = 0;
parameter W34TO3 = 0;
parameter W34TO4 = 0;
parameter W34TO5 = 0;
parameter W34TO6 = 0;
parameter W34TO7 = 0;
parameter W34TO8 = 0;
parameter W34TO9 = 0;
parameter W34TO10 = 0;
parameter W34TO11 = 0;
parameter W34TO12 = 0;
parameter W34TO13 = 0;
parameter W34TO14 = 0;
parameter W34TO15 = 0;
parameter W34TO16 = 0;
parameter W34TO17 = 0;
parameter W34TO18 = 0;
parameter W34TO19 = 0;
parameter W34TO20 = 0;
parameter W34TO21 = 0;
parameter W34TO22 = 0;
parameter W34TO23 = 0;
parameter W34TO24 = 0;
parameter W34TO25 = 0;
parameter W34TO26 = 0;
parameter W34TO27 = 0;
parameter W34TO28 = 0;
parameter W34TO29 = 0;
parameter W34TO30 = 0;
parameter W34TO31 = 0;
parameter W34TO32 = 0;
parameter W34TO33 = 0;
parameter W34TO34 = 0;
parameter W34TO35 = 0;
parameter W34TO36 = 0;
parameter W34TO37 = 0;
parameter W34TO38 = 0;
parameter W34TO39 = 0;
parameter W34TO40 = 0;
parameter W34TO41 = 0;
parameter W34TO42 = 0;
parameter W34TO43 = 0;
parameter W34TO44 = 0;
parameter W34TO45 = 0;
parameter W34TO46 = 0;
parameter W34TO47 = 0;
parameter W34TO48 = 0;
parameter W34TO49 = 0;
parameter W34TO50 = 0;
parameter W34TO51 = 0;
parameter W34TO52 = 0;
parameter W34TO53 = 0;
parameter W34TO54 = 0;
parameter W34TO55 = 0;
parameter W34TO56 = 0;
parameter W34TO57 = 0;
parameter W34TO58 = 0;
parameter W34TO59 = 0;
parameter W34TO60 = 0;
parameter W34TO61 = 0;
parameter W34TO62 = 0;
parameter W34TO63 = 0;
parameter W34TO64 = 0;
parameter W34TO65 = 0;
parameter W34TO66 = 0;
parameter W34TO67 = 0;
parameter W34TO68 = 0;
parameter W34TO69 = 0;
parameter W34TO70 = 0;
parameter W34TO71 = 0;
parameter W34TO72 = 0;
parameter W34TO73 = 0;
parameter W34TO74 = 0;
parameter W34TO75 = 0;
parameter W34TO76 = 0;
parameter W34TO77 = 0;
parameter W34TO78 = 0;
parameter W34TO79 = 0;
parameter W34TO80 = 0;
parameter W34TO81 = 0;
parameter W34TO82 = 0;
parameter W34TO83 = 0;
parameter W34TO84 = 0;
parameter W34TO85 = 0;
parameter W34TO86 = 0;
parameter W34TO87 = 0;
parameter W34TO88 = 0;
parameter W34TO89 = 0;
parameter W34TO90 = 0;
parameter W34TO91 = 0;
parameter W34TO92 = 0;
parameter W34TO93 = 0;
parameter W34TO94 = 0;
parameter W34TO95 = 0;
parameter W34TO96 = 0;
parameter W34TO97 = 0;
parameter W34TO98 = 0;
parameter W34TO99 = 0;
parameter W35TO0 = 0;
parameter W35TO1 = 0;
parameter W35TO2 = 0;
parameter W35TO3 = 0;
parameter W35TO4 = 0;
parameter W35TO5 = 0;
parameter W35TO6 = 0;
parameter W35TO7 = 0;
parameter W35TO8 = 0;
parameter W35TO9 = 0;
parameter W35TO10 = 0;
parameter W35TO11 = 0;
parameter W35TO12 = 0;
parameter W35TO13 = 0;
parameter W35TO14 = 0;
parameter W35TO15 = 0;
parameter W35TO16 = 0;
parameter W35TO17 = 0;
parameter W35TO18 = 0;
parameter W35TO19 = 0;
parameter W35TO20 = 0;
parameter W35TO21 = 0;
parameter W35TO22 = 0;
parameter W35TO23 = 0;
parameter W35TO24 = 0;
parameter W35TO25 = 0;
parameter W35TO26 = 0;
parameter W35TO27 = 0;
parameter W35TO28 = 0;
parameter W35TO29 = 0;
parameter W35TO30 = 0;
parameter W35TO31 = 0;
parameter W35TO32 = 0;
parameter W35TO33 = 0;
parameter W35TO34 = 0;
parameter W35TO35 = 0;
parameter W35TO36 = 0;
parameter W35TO37 = 0;
parameter W35TO38 = 0;
parameter W35TO39 = 0;
parameter W35TO40 = 0;
parameter W35TO41 = 0;
parameter W35TO42 = 0;
parameter W35TO43 = 0;
parameter W35TO44 = 0;
parameter W35TO45 = 0;
parameter W35TO46 = 0;
parameter W35TO47 = 0;
parameter W35TO48 = 0;
parameter W35TO49 = 0;
parameter W35TO50 = 0;
parameter W35TO51 = 0;
parameter W35TO52 = 0;
parameter W35TO53 = 0;
parameter W35TO54 = 0;
parameter W35TO55 = 0;
parameter W35TO56 = 0;
parameter W35TO57 = 0;
parameter W35TO58 = 0;
parameter W35TO59 = 0;
parameter W35TO60 = 0;
parameter W35TO61 = 0;
parameter W35TO62 = 0;
parameter W35TO63 = 0;
parameter W35TO64 = 0;
parameter W35TO65 = 0;
parameter W35TO66 = 0;
parameter W35TO67 = 0;
parameter W35TO68 = 0;
parameter W35TO69 = 0;
parameter W35TO70 = 0;
parameter W35TO71 = 0;
parameter W35TO72 = 0;
parameter W35TO73 = 0;
parameter W35TO74 = 0;
parameter W35TO75 = 0;
parameter W35TO76 = 0;
parameter W35TO77 = 0;
parameter W35TO78 = 0;
parameter W35TO79 = 0;
parameter W35TO80 = 0;
parameter W35TO81 = 0;
parameter W35TO82 = 0;
parameter W35TO83 = 0;
parameter W35TO84 = 0;
parameter W35TO85 = 0;
parameter W35TO86 = 0;
parameter W35TO87 = 0;
parameter W35TO88 = 0;
parameter W35TO89 = 0;
parameter W35TO90 = 0;
parameter W35TO91 = 0;
parameter W35TO92 = 0;
parameter W35TO93 = 0;
parameter W35TO94 = 0;
parameter W35TO95 = 0;
parameter W35TO96 = 0;
parameter W35TO97 = 0;
parameter W35TO98 = 0;
parameter W35TO99 = 0;
parameter W36TO0 = 0;
parameter W36TO1 = 0;
parameter W36TO2 = 0;
parameter W36TO3 = 0;
parameter W36TO4 = 0;
parameter W36TO5 = 0;
parameter W36TO6 = 0;
parameter W36TO7 = 0;
parameter W36TO8 = 0;
parameter W36TO9 = 0;
parameter W36TO10 = 0;
parameter W36TO11 = 0;
parameter W36TO12 = 0;
parameter W36TO13 = 0;
parameter W36TO14 = 0;
parameter W36TO15 = 0;
parameter W36TO16 = 0;
parameter W36TO17 = 0;
parameter W36TO18 = 0;
parameter W36TO19 = 0;
parameter W36TO20 = 0;
parameter W36TO21 = 0;
parameter W36TO22 = 0;
parameter W36TO23 = 0;
parameter W36TO24 = 0;
parameter W36TO25 = 0;
parameter W36TO26 = 0;
parameter W36TO27 = 0;
parameter W36TO28 = 0;
parameter W36TO29 = 0;
parameter W36TO30 = 0;
parameter W36TO31 = 0;
parameter W36TO32 = 0;
parameter W36TO33 = 0;
parameter W36TO34 = 0;
parameter W36TO35 = 0;
parameter W36TO36 = 0;
parameter W36TO37 = 0;
parameter W36TO38 = 0;
parameter W36TO39 = 0;
parameter W36TO40 = 0;
parameter W36TO41 = 0;
parameter W36TO42 = 0;
parameter W36TO43 = 0;
parameter W36TO44 = 0;
parameter W36TO45 = 0;
parameter W36TO46 = 0;
parameter W36TO47 = 0;
parameter W36TO48 = 0;
parameter W36TO49 = 0;
parameter W36TO50 = 0;
parameter W36TO51 = 0;
parameter W36TO52 = 0;
parameter W36TO53 = 0;
parameter W36TO54 = 0;
parameter W36TO55 = 0;
parameter W36TO56 = 0;
parameter W36TO57 = 0;
parameter W36TO58 = 0;
parameter W36TO59 = 0;
parameter W36TO60 = 0;
parameter W36TO61 = 0;
parameter W36TO62 = 0;
parameter W36TO63 = 0;
parameter W36TO64 = 0;
parameter W36TO65 = 0;
parameter W36TO66 = 0;
parameter W36TO67 = 0;
parameter W36TO68 = 0;
parameter W36TO69 = 0;
parameter W36TO70 = 0;
parameter W36TO71 = 0;
parameter W36TO72 = 0;
parameter W36TO73 = 0;
parameter W36TO74 = 0;
parameter W36TO75 = 0;
parameter W36TO76 = 0;
parameter W36TO77 = 0;
parameter W36TO78 = 0;
parameter W36TO79 = 0;
parameter W36TO80 = 0;
parameter W36TO81 = 0;
parameter W36TO82 = 0;
parameter W36TO83 = 0;
parameter W36TO84 = 0;
parameter W36TO85 = 0;
parameter W36TO86 = 0;
parameter W36TO87 = 0;
parameter W36TO88 = 0;
parameter W36TO89 = 0;
parameter W36TO90 = 0;
parameter W36TO91 = 0;
parameter W36TO92 = 0;
parameter W36TO93 = 0;
parameter W36TO94 = 0;
parameter W36TO95 = 0;
parameter W36TO96 = 0;
parameter W36TO97 = 0;
parameter W36TO98 = 0;
parameter W36TO99 = 0;
parameter W37TO0 = 0;
parameter W37TO1 = 0;
parameter W37TO2 = 0;
parameter W37TO3 = 0;
parameter W37TO4 = 0;
parameter W37TO5 = 0;
parameter W37TO6 = 0;
parameter W37TO7 = 0;
parameter W37TO8 = 0;
parameter W37TO9 = 0;
parameter W37TO10 = 0;
parameter W37TO11 = 0;
parameter W37TO12 = 0;
parameter W37TO13 = 0;
parameter W37TO14 = 0;
parameter W37TO15 = 0;
parameter W37TO16 = 0;
parameter W37TO17 = 0;
parameter W37TO18 = 0;
parameter W37TO19 = 0;
parameter W37TO20 = 0;
parameter W37TO21 = 0;
parameter W37TO22 = 0;
parameter W37TO23 = 0;
parameter W37TO24 = 0;
parameter W37TO25 = 0;
parameter W37TO26 = 0;
parameter W37TO27 = 0;
parameter W37TO28 = 0;
parameter W37TO29 = 0;
parameter W37TO30 = 0;
parameter W37TO31 = 0;
parameter W37TO32 = 0;
parameter W37TO33 = 0;
parameter W37TO34 = 0;
parameter W37TO35 = 0;
parameter W37TO36 = 0;
parameter W37TO37 = 0;
parameter W37TO38 = 0;
parameter W37TO39 = 0;
parameter W37TO40 = 0;
parameter W37TO41 = 0;
parameter W37TO42 = 0;
parameter W37TO43 = 0;
parameter W37TO44 = 0;
parameter W37TO45 = 0;
parameter W37TO46 = 0;
parameter W37TO47 = 0;
parameter W37TO48 = 0;
parameter W37TO49 = 0;
parameter W37TO50 = 0;
parameter W37TO51 = 0;
parameter W37TO52 = 0;
parameter W37TO53 = 0;
parameter W37TO54 = 0;
parameter W37TO55 = 0;
parameter W37TO56 = 0;
parameter W37TO57 = 0;
parameter W37TO58 = 0;
parameter W37TO59 = 0;
parameter W37TO60 = 0;
parameter W37TO61 = 0;
parameter W37TO62 = 0;
parameter W37TO63 = 0;
parameter W37TO64 = 0;
parameter W37TO65 = 0;
parameter W37TO66 = 0;
parameter W37TO67 = 0;
parameter W37TO68 = 0;
parameter W37TO69 = 0;
parameter W37TO70 = 0;
parameter W37TO71 = 0;
parameter W37TO72 = 0;
parameter W37TO73 = 0;
parameter W37TO74 = 0;
parameter W37TO75 = 0;
parameter W37TO76 = 0;
parameter W37TO77 = 0;
parameter W37TO78 = 0;
parameter W37TO79 = 0;
parameter W37TO80 = 0;
parameter W37TO81 = 0;
parameter W37TO82 = 0;
parameter W37TO83 = 0;
parameter W37TO84 = 0;
parameter W37TO85 = 0;
parameter W37TO86 = 0;
parameter W37TO87 = 0;
parameter W37TO88 = 0;
parameter W37TO89 = 0;
parameter W37TO90 = 0;
parameter W37TO91 = 0;
parameter W37TO92 = 0;
parameter W37TO93 = 0;
parameter W37TO94 = 0;
parameter W37TO95 = 0;
parameter W37TO96 = 0;
parameter W37TO97 = 0;
parameter W37TO98 = 0;
parameter W37TO99 = 0;
parameter W38TO0 = 0;
parameter W38TO1 = 0;
parameter W38TO2 = 0;
parameter W38TO3 = 0;
parameter W38TO4 = 0;
parameter W38TO5 = 0;
parameter W38TO6 = 0;
parameter W38TO7 = 0;
parameter W38TO8 = 0;
parameter W38TO9 = 0;
parameter W38TO10 = 0;
parameter W38TO11 = 0;
parameter W38TO12 = 0;
parameter W38TO13 = 0;
parameter W38TO14 = 0;
parameter W38TO15 = 0;
parameter W38TO16 = 0;
parameter W38TO17 = 0;
parameter W38TO18 = 0;
parameter W38TO19 = 0;
parameter W38TO20 = 0;
parameter W38TO21 = 0;
parameter W38TO22 = 0;
parameter W38TO23 = 0;
parameter W38TO24 = 0;
parameter W38TO25 = 0;
parameter W38TO26 = 0;
parameter W38TO27 = 0;
parameter W38TO28 = 0;
parameter W38TO29 = 0;
parameter W38TO30 = 0;
parameter W38TO31 = 0;
parameter W38TO32 = 0;
parameter W38TO33 = 0;
parameter W38TO34 = 0;
parameter W38TO35 = 0;
parameter W38TO36 = 0;
parameter W38TO37 = 0;
parameter W38TO38 = 0;
parameter W38TO39 = 0;
parameter W38TO40 = 0;
parameter W38TO41 = 0;
parameter W38TO42 = 0;
parameter W38TO43 = 0;
parameter W38TO44 = 0;
parameter W38TO45 = 0;
parameter W38TO46 = 0;
parameter W38TO47 = 0;
parameter W38TO48 = 0;
parameter W38TO49 = 0;
parameter W38TO50 = 0;
parameter W38TO51 = 0;
parameter W38TO52 = 0;
parameter W38TO53 = 0;
parameter W38TO54 = 0;
parameter W38TO55 = 0;
parameter W38TO56 = 0;
parameter W38TO57 = 0;
parameter W38TO58 = 0;
parameter W38TO59 = 0;
parameter W38TO60 = 0;
parameter W38TO61 = 0;
parameter W38TO62 = 0;
parameter W38TO63 = 0;
parameter W38TO64 = 0;
parameter W38TO65 = 0;
parameter W38TO66 = 0;
parameter W38TO67 = 0;
parameter W38TO68 = 0;
parameter W38TO69 = 0;
parameter W38TO70 = 0;
parameter W38TO71 = 0;
parameter W38TO72 = 0;
parameter W38TO73 = 0;
parameter W38TO74 = 0;
parameter W38TO75 = 0;
parameter W38TO76 = 0;
parameter W38TO77 = 0;
parameter W38TO78 = 0;
parameter W38TO79 = 0;
parameter W38TO80 = 0;
parameter W38TO81 = 0;
parameter W38TO82 = 0;
parameter W38TO83 = 0;
parameter W38TO84 = 0;
parameter W38TO85 = 0;
parameter W38TO86 = 0;
parameter W38TO87 = 0;
parameter W38TO88 = 0;
parameter W38TO89 = 0;
parameter W38TO90 = 0;
parameter W38TO91 = 0;
parameter W38TO92 = 0;
parameter W38TO93 = 0;
parameter W38TO94 = 0;
parameter W38TO95 = 0;
parameter W38TO96 = 0;
parameter W38TO97 = 0;
parameter W38TO98 = 0;
parameter W38TO99 = 0;
parameter W39TO0 = 0;
parameter W39TO1 = 0;
parameter W39TO2 = 0;
parameter W39TO3 = 0;
parameter W39TO4 = 0;
parameter W39TO5 = 0;
parameter W39TO6 = 0;
parameter W39TO7 = 0;
parameter W39TO8 = 0;
parameter W39TO9 = 0;
parameter W39TO10 = 0;
parameter W39TO11 = 0;
parameter W39TO12 = 0;
parameter W39TO13 = 0;
parameter W39TO14 = 0;
parameter W39TO15 = 0;
parameter W39TO16 = 0;
parameter W39TO17 = 0;
parameter W39TO18 = 0;
parameter W39TO19 = 0;
parameter W39TO20 = 0;
parameter W39TO21 = 0;
parameter W39TO22 = 0;
parameter W39TO23 = 0;
parameter W39TO24 = 0;
parameter W39TO25 = 0;
parameter W39TO26 = 0;
parameter W39TO27 = 0;
parameter W39TO28 = 0;
parameter W39TO29 = 0;
parameter W39TO30 = 0;
parameter W39TO31 = 0;
parameter W39TO32 = 0;
parameter W39TO33 = 0;
parameter W39TO34 = 0;
parameter W39TO35 = 0;
parameter W39TO36 = 0;
parameter W39TO37 = 0;
parameter W39TO38 = 0;
parameter W39TO39 = 0;
parameter W39TO40 = 0;
parameter W39TO41 = 0;
parameter W39TO42 = 0;
parameter W39TO43 = 0;
parameter W39TO44 = 0;
parameter W39TO45 = 0;
parameter W39TO46 = 0;
parameter W39TO47 = 0;
parameter W39TO48 = 0;
parameter W39TO49 = 0;
parameter W39TO50 = 0;
parameter W39TO51 = 0;
parameter W39TO52 = 0;
parameter W39TO53 = 0;
parameter W39TO54 = 0;
parameter W39TO55 = 0;
parameter W39TO56 = 0;
parameter W39TO57 = 0;
parameter W39TO58 = 0;
parameter W39TO59 = 0;
parameter W39TO60 = 0;
parameter W39TO61 = 0;
parameter W39TO62 = 0;
parameter W39TO63 = 0;
parameter W39TO64 = 0;
parameter W39TO65 = 0;
parameter W39TO66 = 0;
parameter W39TO67 = 0;
parameter W39TO68 = 0;
parameter W39TO69 = 0;
parameter W39TO70 = 0;
parameter W39TO71 = 0;
parameter W39TO72 = 0;
parameter W39TO73 = 0;
parameter W39TO74 = 0;
parameter W39TO75 = 0;
parameter W39TO76 = 0;
parameter W39TO77 = 0;
parameter W39TO78 = 0;
parameter W39TO79 = 0;
parameter W39TO80 = 0;
parameter W39TO81 = 0;
parameter W39TO82 = 0;
parameter W39TO83 = 0;
parameter W39TO84 = 0;
parameter W39TO85 = 0;
parameter W39TO86 = 0;
parameter W39TO87 = 0;
parameter W39TO88 = 0;
parameter W39TO89 = 0;
parameter W39TO90 = 0;
parameter W39TO91 = 0;
parameter W39TO92 = 0;
parameter W39TO93 = 0;
parameter W39TO94 = 0;
parameter W39TO95 = 0;
parameter W39TO96 = 0;
parameter W39TO97 = 0;
parameter W39TO98 = 0;
parameter W39TO99 = 0;
parameter W40TO0 = 0;
parameter W40TO1 = 0;
parameter W40TO2 = 0;
parameter W40TO3 = 0;
parameter W40TO4 = 0;
parameter W40TO5 = 0;
parameter W40TO6 = 0;
parameter W40TO7 = 0;
parameter W40TO8 = 0;
parameter W40TO9 = 0;
parameter W40TO10 = 0;
parameter W40TO11 = 0;
parameter W40TO12 = 0;
parameter W40TO13 = 0;
parameter W40TO14 = 0;
parameter W40TO15 = 0;
parameter W40TO16 = 0;
parameter W40TO17 = 0;
parameter W40TO18 = 0;
parameter W40TO19 = 0;
parameter W40TO20 = 0;
parameter W40TO21 = 0;
parameter W40TO22 = 0;
parameter W40TO23 = 0;
parameter W40TO24 = 0;
parameter W40TO25 = 0;
parameter W40TO26 = 0;
parameter W40TO27 = 0;
parameter W40TO28 = 0;
parameter W40TO29 = 0;
parameter W40TO30 = 0;
parameter W40TO31 = 0;
parameter W40TO32 = 0;
parameter W40TO33 = 0;
parameter W40TO34 = 0;
parameter W40TO35 = 0;
parameter W40TO36 = 0;
parameter W40TO37 = 0;
parameter W40TO38 = 0;
parameter W40TO39 = 0;
parameter W40TO40 = 0;
parameter W40TO41 = 0;
parameter W40TO42 = 0;
parameter W40TO43 = 0;
parameter W40TO44 = 0;
parameter W40TO45 = 0;
parameter W40TO46 = 0;
parameter W40TO47 = 0;
parameter W40TO48 = 0;
parameter W40TO49 = 0;
parameter W40TO50 = 0;
parameter W40TO51 = 0;
parameter W40TO52 = 0;
parameter W40TO53 = 0;
parameter W40TO54 = 0;
parameter W40TO55 = 0;
parameter W40TO56 = 0;
parameter W40TO57 = 0;
parameter W40TO58 = 0;
parameter W40TO59 = 0;
parameter W40TO60 = 0;
parameter W40TO61 = 0;
parameter W40TO62 = 0;
parameter W40TO63 = 0;
parameter W40TO64 = 0;
parameter W40TO65 = 0;
parameter W40TO66 = 0;
parameter W40TO67 = 0;
parameter W40TO68 = 0;
parameter W40TO69 = 0;
parameter W40TO70 = 0;
parameter W40TO71 = 0;
parameter W40TO72 = 0;
parameter W40TO73 = 0;
parameter W40TO74 = 0;
parameter W40TO75 = 0;
parameter W40TO76 = 0;
parameter W40TO77 = 0;
parameter W40TO78 = 0;
parameter W40TO79 = 0;
parameter W40TO80 = 0;
parameter W40TO81 = 0;
parameter W40TO82 = 0;
parameter W40TO83 = 0;
parameter W40TO84 = 0;
parameter W40TO85 = 0;
parameter W40TO86 = 0;
parameter W40TO87 = 0;
parameter W40TO88 = 0;
parameter W40TO89 = 0;
parameter W40TO90 = 0;
parameter W40TO91 = 0;
parameter W40TO92 = 0;
parameter W40TO93 = 0;
parameter W40TO94 = 0;
parameter W40TO95 = 0;
parameter W40TO96 = 0;
parameter W40TO97 = 0;
parameter W40TO98 = 0;
parameter W40TO99 = 0;
parameter W41TO0 = 0;
parameter W41TO1 = 0;
parameter W41TO2 = 0;
parameter W41TO3 = 0;
parameter W41TO4 = 0;
parameter W41TO5 = 0;
parameter W41TO6 = 0;
parameter W41TO7 = 0;
parameter W41TO8 = 0;
parameter W41TO9 = 0;
parameter W41TO10 = 0;
parameter W41TO11 = 0;
parameter W41TO12 = 0;
parameter W41TO13 = 0;
parameter W41TO14 = 0;
parameter W41TO15 = 0;
parameter W41TO16 = 0;
parameter W41TO17 = 0;
parameter W41TO18 = 0;
parameter W41TO19 = 0;
parameter W41TO20 = 0;
parameter W41TO21 = 0;
parameter W41TO22 = 0;
parameter W41TO23 = 0;
parameter W41TO24 = 0;
parameter W41TO25 = 0;
parameter W41TO26 = 0;
parameter W41TO27 = 0;
parameter W41TO28 = 0;
parameter W41TO29 = 0;
parameter W41TO30 = 0;
parameter W41TO31 = 0;
parameter W41TO32 = 0;
parameter W41TO33 = 0;
parameter W41TO34 = 0;
parameter W41TO35 = 0;
parameter W41TO36 = 0;
parameter W41TO37 = 0;
parameter W41TO38 = 0;
parameter W41TO39 = 0;
parameter W41TO40 = 0;
parameter W41TO41 = 0;
parameter W41TO42 = 0;
parameter W41TO43 = 0;
parameter W41TO44 = 0;
parameter W41TO45 = 0;
parameter W41TO46 = 0;
parameter W41TO47 = 0;
parameter W41TO48 = 0;
parameter W41TO49 = 0;
parameter W41TO50 = 0;
parameter W41TO51 = 0;
parameter W41TO52 = 0;
parameter W41TO53 = 0;
parameter W41TO54 = 0;
parameter W41TO55 = 0;
parameter W41TO56 = 0;
parameter W41TO57 = 0;
parameter W41TO58 = 0;
parameter W41TO59 = 0;
parameter W41TO60 = 0;
parameter W41TO61 = 0;
parameter W41TO62 = 0;
parameter W41TO63 = 0;
parameter W41TO64 = 0;
parameter W41TO65 = 0;
parameter W41TO66 = 0;
parameter W41TO67 = 0;
parameter W41TO68 = 0;
parameter W41TO69 = 0;
parameter W41TO70 = 0;
parameter W41TO71 = 0;
parameter W41TO72 = 0;
parameter W41TO73 = 0;
parameter W41TO74 = 0;
parameter W41TO75 = 0;
parameter W41TO76 = 0;
parameter W41TO77 = 0;
parameter W41TO78 = 0;
parameter W41TO79 = 0;
parameter W41TO80 = 0;
parameter W41TO81 = 0;
parameter W41TO82 = 0;
parameter W41TO83 = 0;
parameter W41TO84 = 0;
parameter W41TO85 = 0;
parameter W41TO86 = 0;
parameter W41TO87 = 0;
parameter W41TO88 = 0;
parameter W41TO89 = 0;
parameter W41TO90 = 0;
parameter W41TO91 = 0;
parameter W41TO92 = 0;
parameter W41TO93 = 0;
parameter W41TO94 = 0;
parameter W41TO95 = 0;
parameter W41TO96 = 0;
parameter W41TO97 = 0;
parameter W41TO98 = 0;
parameter W41TO99 = 0;
parameter W42TO0 = 0;
parameter W42TO1 = 0;
parameter W42TO2 = 0;
parameter W42TO3 = 0;
parameter W42TO4 = 0;
parameter W42TO5 = 0;
parameter W42TO6 = 0;
parameter W42TO7 = 0;
parameter W42TO8 = 0;
parameter W42TO9 = 0;
parameter W42TO10 = 0;
parameter W42TO11 = 0;
parameter W42TO12 = 0;
parameter W42TO13 = 0;
parameter W42TO14 = 0;
parameter W42TO15 = 0;
parameter W42TO16 = 0;
parameter W42TO17 = 0;
parameter W42TO18 = 0;
parameter W42TO19 = 0;
parameter W42TO20 = 0;
parameter W42TO21 = 0;
parameter W42TO22 = 0;
parameter W42TO23 = 0;
parameter W42TO24 = 0;
parameter W42TO25 = 0;
parameter W42TO26 = 0;
parameter W42TO27 = 0;
parameter W42TO28 = 0;
parameter W42TO29 = 0;
parameter W42TO30 = 0;
parameter W42TO31 = 0;
parameter W42TO32 = 0;
parameter W42TO33 = 0;
parameter W42TO34 = 0;
parameter W42TO35 = 0;
parameter W42TO36 = 0;
parameter W42TO37 = 0;
parameter W42TO38 = 0;
parameter W42TO39 = 0;
parameter W42TO40 = 0;
parameter W42TO41 = 0;
parameter W42TO42 = 0;
parameter W42TO43 = 0;
parameter W42TO44 = 0;
parameter W42TO45 = 0;
parameter W42TO46 = 0;
parameter W42TO47 = 0;
parameter W42TO48 = 0;
parameter W42TO49 = 0;
parameter W42TO50 = 0;
parameter W42TO51 = 0;
parameter W42TO52 = 0;
parameter W42TO53 = 0;
parameter W42TO54 = 0;
parameter W42TO55 = 0;
parameter W42TO56 = 0;
parameter W42TO57 = 0;
parameter W42TO58 = 0;
parameter W42TO59 = 0;
parameter W42TO60 = 0;
parameter W42TO61 = 0;
parameter W42TO62 = 0;
parameter W42TO63 = 0;
parameter W42TO64 = 0;
parameter W42TO65 = 0;
parameter W42TO66 = 0;
parameter W42TO67 = 0;
parameter W42TO68 = 0;
parameter W42TO69 = 0;
parameter W42TO70 = 0;
parameter W42TO71 = 0;
parameter W42TO72 = 0;
parameter W42TO73 = 0;
parameter W42TO74 = 0;
parameter W42TO75 = 0;
parameter W42TO76 = 0;
parameter W42TO77 = 0;
parameter W42TO78 = 0;
parameter W42TO79 = 0;
parameter W42TO80 = 0;
parameter W42TO81 = 0;
parameter W42TO82 = 0;
parameter W42TO83 = 0;
parameter W42TO84 = 0;
parameter W42TO85 = 0;
parameter W42TO86 = 0;
parameter W42TO87 = 0;
parameter W42TO88 = 0;
parameter W42TO89 = 0;
parameter W42TO90 = 0;
parameter W42TO91 = 0;
parameter W42TO92 = 0;
parameter W42TO93 = 0;
parameter W42TO94 = 0;
parameter W42TO95 = 0;
parameter W42TO96 = 0;
parameter W42TO97 = 0;
parameter W42TO98 = 0;
parameter W42TO99 = 0;
parameter W43TO0 = 0;
parameter W43TO1 = 0;
parameter W43TO2 = 0;
parameter W43TO3 = 0;
parameter W43TO4 = 0;
parameter W43TO5 = 0;
parameter W43TO6 = 0;
parameter W43TO7 = 0;
parameter W43TO8 = 0;
parameter W43TO9 = 0;
parameter W43TO10 = 0;
parameter W43TO11 = 0;
parameter W43TO12 = 0;
parameter W43TO13 = 0;
parameter W43TO14 = 0;
parameter W43TO15 = 0;
parameter W43TO16 = 0;
parameter W43TO17 = 0;
parameter W43TO18 = 0;
parameter W43TO19 = 0;
parameter W43TO20 = 0;
parameter W43TO21 = 0;
parameter W43TO22 = 0;
parameter W43TO23 = 0;
parameter W43TO24 = 0;
parameter W43TO25 = 0;
parameter W43TO26 = 0;
parameter W43TO27 = 0;
parameter W43TO28 = 0;
parameter W43TO29 = 0;
parameter W43TO30 = 0;
parameter W43TO31 = 0;
parameter W43TO32 = 0;
parameter W43TO33 = 0;
parameter W43TO34 = 0;
parameter W43TO35 = 0;
parameter W43TO36 = 0;
parameter W43TO37 = 0;
parameter W43TO38 = 0;
parameter W43TO39 = 0;
parameter W43TO40 = 0;
parameter W43TO41 = 0;
parameter W43TO42 = 0;
parameter W43TO43 = 0;
parameter W43TO44 = 0;
parameter W43TO45 = 0;
parameter W43TO46 = 0;
parameter W43TO47 = 0;
parameter W43TO48 = 0;
parameter W43TO49 = 0;
parameter W43TO50 = 0;
parameter W43TO51 = 0;
parameter W43TO52 = 0;
parameter W43TO53 = 0;
parameter W43TO54 = 0;
parameter W43TO55 = 0;
parameter W43TO56 = 0;
parameter W43TO57 = 0;
parameter W43TO58 = 0;
parameter W43TO59 = 0;
parameter W43TO60 = 0;
parameter W43TO61 = 0;
parameter W43TO62 = 0;
parameter W43TO63 = 0;
parameter W43TO64 = 0;
parameter W43TO65 = 0;
parameter W43TO66 = 0;
parameter W43TO67 = 0;
parameter W43TO68 = 0;
parameter W43TO69 = 0;
parameter W43TO70 = 0;
parameter W43TO71 = 0;
parameter W43TO72 = 0;
parameter W43TO73 = 0;
parameter W43TO74 = 0;
parameter W43TO75 = 0;
parameter W43TO76 = 0;
parameter W43TO77 = 0;
parameter W43TO78 = 0;
parameter W43TO79 = 0;
parameter W43TO80 = 0;
parameter W43TO81 = 0;
parameter W43TO82 = 0;
parameter W43TO83 = 0;
parameter W43TO84 = 0;
parameter W43TO85 = 0;
parameter W43TO86 = 0;
parameter W43TO87 = 0;
parameter W43TO88 = 0;
parameter W43TO89 = 0;
parameter W43TO90 = 0;
parameter W43TO91 = 0;
parameter W43TO92 = 0;
parameter W43TO93 = 0;
parameter W43TO94 = 0;
parameter W43TO95 = 0;
parameter W43TO96 = 0;
parameter W43TO97 = 0;
parameter W43TO98 = 0;
parameter W43TO99 = 0;
parameter W44TO0 = 0;
parameter W44TO1 = 0;
parameter W44TO2 = 0;
parameter W44TO3 = 0;
parameter W44TO4 = 0;
parameter W44TO5 = 0;
parameter W44TO6 = 0;
parameter W44TO7 = 0;
parameter W44TO8 = 0;
parameter W44TO9 = 0;
parameter W44TO10 = 0;
parameter W44TO11 = 0;
parameter W44TO12 = 0;
parameter W44TO13 = 0;
parameter W44TO14 = 0;
parameter W44TO15 = 0;
parameter W44TO16 = 0;
parameter W44TO17 = 0;
parameter W44TO18 = 0;
parameter W44TO19 = 0;
parameter W44TO20 = 0;
parameter W44TO21 = 0;
parameter W44TO22 = 0;
parameter W44TO23 = 0;
parameter W44TO24 = 0;
parameter W44TO25 = 0;
parameter W44TO26 = 0;
parameter W44TO27 = 0;
parameter W44TO28 = 0;
parameter W44TO29 = 0;
parameter W44TO30 = 0;
parameter W44TO31 = 0;
parameter W44TO32 = 0;
parameter W44TO33 = 0;
parameter W44TO34 = 0;
parameter W44TO35 = 0;
parameter W44TO36 = 0;
parameter W44TO37 = 0;
parameter W44TO38 = 0;
parameter W44TO39 = 0;
parameter W44TO40 = 0;
parameter W44TO41 = 0;
parameter W44TO42 = 0;
parameter W44TO43 = 0;
parameter W44TO44 = 0;
parameter W44TO45 = 0;
parameter W44TO46 = 0;
parameter W44TO47 = 0;
parameter W44TO48 = 0;
parameter W44TO49 = 0;
parameter W44TO50 = 0;
parameter W44TO51 = 0;
parameter W44TO52 = 0;
parameter W44TO53 = 0;
parameter W44TO54 = 0;
parameter W44TO55 = 0;
parameter W44TO56 = 0;
parameter W44TO57 = 0;
parameter W44TO58 = 0;
parameter W44TO59 = 0;
parameter W44TO60 = 0;
parameter W44TO61 = 0;
parameter W44TO62 = 0;
parameter W44TO63 = 0;
parameter W44TO64 = 0;
parameter W44TO65 = 0;
parameter W44TO66 = 0;
parameter W44TO67 = 0;
parameter W44TO68 = 0;
parameter W44TO69 = 0;
parameter W44TO70 = 0;
parameter W44TO71 = 0;
parameter W44TO72 = 0;
parameter W44TO73 = 0;
parameter W44TO74 = 0;
parameter W44TO75 = 0;
parameter W44TO76 = 0;
parameter W44TO77 = 0;
parameter W44TO78 = 0;
parameter W44TO79 = 0;
parameter W44TO80 = 0;
parameter W44TO81 = 0;
parameter W44TO82 = 0;
parameter W44TO83 = 0;
parameter W44TO84 = 0;
parameter W44TO85 = 0;
parameter W44TO86 = 0;
parameter W44TO87 = 0;
parameter W44TO88 = 0;
parameter W44TO89 = 0;
parameter W44TO90 = 0;
parameter W44TO91 = 0;
parameter W44TO92 = 0;
parameter W44TO93 = 0;
parameter W44TO94 = 0;
parameter W44TO95 = 0;
parameter W44TO96 = 0;
parameter W44TO97 = 0;
parameter W44TO98 = 0;
parameter W44TO99 = 0;
parameter W45TO0 = 0;
parameter W45TO1 = 0;
parameter W45TO2 = 0;
parameter W45TO3 = 0;
parameter W45TO4 = 0;
parameter W45TO5 = 0;
parameter W45TO6 = 0;
parameter W45TO7 = 0;
parameter W45TO8 = 0;
parameter W45TO9 = 0;
parameter W45TO10 = 0;
parameter W45TO11 = 0;
parameter W45TO12 = 0;
parameter W45TO13 = 0;
parameter W45TO14 = 0;
parameter W45TO15 = 0;
parameter W45TO16 = 0;
parameter W45TO17 = 0;
parameter W45TO18 = 0;
parameter W45TO19 = 0;
parameter W45TO20 = 0;
parameter W45TO21 = 0;
parameter W45TO22 = 0;
parameter W45TO23 = 0;
parameter W45TO24 = 0;
parameter W45TO25 = 0;
parameter W45TO26 = 0;
parameter W45TO27 = 0;
parameter W45TO28 = 0;
parameter W45TO29 = 0;
parameter W45TO30 = 0;
parameter W45TO31 = 0;
parameter W45TO32 = 0;
parameter W45TO33 = 0;
parameter W45TO34 = 0;
parameter W45TO35 = 0;
parameter W45TO36 = 0;
parameter W45TO37 = 0;
parameter W45TO38 = 0;
parameter W45TO39 = 0;
parameter W45TO40 = 0;
parameter W45TO41 = 0;
parameter W45TO42 = 0;
parameter W45TO43 = 0;
parameter W45TO44 = 0;
parameter W45TO45 = 0;
parameter W45TO46 = 0;
parameter W45TO47 = 0;
parameter W45TO48 = 0;
parameter W45TO49 = 0;
parameter W45TO50 = 0;
parameter W45TO51 = 0;
parameter W45TO52 = 0;
parameter W45TO53 = 0;
parameter W45TO54 = 0;
parameter W45TO55 = 0;
parameter W45TO56 = 0;
parameter W45TO57 = 0;
parameter W45TO58 = 0;
parameter W45TO59 = 0;
parameter W45TO60 = 0;
parameter W45TO61 = 0;
parameter W45TO62 = 0;
parameter W45TO63 = 0;
parameter W45TO64 = 0;
parameter W45TO65 = 0;
parameter W45TO66 = 0;
parameter W45TO67 = 0;
parameter W45TO68 = 0;
parameter W45TO69 = 0;
parameter W45TO70 = 0;
parameter W45TO71 = 0;
parameter W45TO72 = 0;
parameter W45TO73 = 0;
parameter W45TO74 = 0;
parameter W45TO75 = 0;
parameter W45TO76 = 0;
parameter W45TO77 = 0;
parameter W45TO78 = 0;
parameter W45TO79 = 0;
parameter W45TO80 = 0;
parameter W45TO81 = 0;
parameter W45TO82 = 0;
parameter W45TO83 = 0;
parameter W45TO84 = 0;
parameter W45TO85 = 0;
parameter W45TO86 = 0;
parameter W45TO87 = 0;
parameter W45TO88 = 0;
parameter W45TO89 = 0;
parameter W45TO90 = 0;
parameter W45TO91 = 0;
parameter W45TO92 = 0;
parameter W45TO93 = 0;
parameter W45TO94 = 0;
parameter W45TO95 = 0;
parameter W45TO96 = 0;
parameter W45TO97 = 0;
parameter W45TO98 = 0;
parameter W45TO99 = 0;
parameter W46TO0 = 0;
parameter W46TO1 = 0;
parameter W46TO2 = 0;
parameter W46TO3 = 0;
parameter W46TO4 = 0;
parameter W46TO5 = 0;
parameter W46TO6 = 0;
parameter W46TO7 = 0;
parameter W46TO8 = 0;
parameter W46TO9 = 0;
parameter W46TO10 = 0;
parameter W46TO11 = 0;
parameter W46TO12 = 0;
parameter W46TO13 = 0;
parameter W46TO14 = 0;
parameter W46TO15 = 0;
parameter W46TO16 = 0;
parameter W46TO17 = 0;
parameter W46TO18 = 0;
parameter W46TO19 = 0;
parameter W46TO20 = 0;
parameter W46TO21 = 0;
parameter W46TO22 = 0;
parameter W46TO23 = 0;
parameter W46TO24 = 0;
parameter W46TO25 = 0;
parameter W46TO26 = 0;
parameter W46TO27 = 0;
parameter W46TO28 = 0;
parameter W46TO29 = 0;
parameter W46TO30 = 0;
parameter W46TO31 = 0;
parameter W46TO32 = 0;
parameter W46TO33 = 0;
parameter W46TO34 = 0;
parameter W46TO35 = 0;
parameter W46TO36 = 0;
parameter W46TO37 = 0;
parameter W46TO38 = 0;
parameter W46TO39 = 0;
parameter W46TO40 = 0;
parameter W46TO41 = 0;
parameter W46TO42 = 0;
parameter W46TO43 = 0;
parameter W46TO44 = 0;
parameter W46TO45 = 0;
parameter W46TO46 = 0;
parameter W46TO47 = 0;
parameter W46TO48 = 0;
parameter W46TO49 = 0;
parameter W46TO50 = 0;
parameter W46TO51 = 0;
parameter W46TO52 = 0;
parameter W46TO53 = 0;
parameter W46TO54 = 0;
parameter W46TO55 = 0;
parameter W46TO56 = 0;
parameter W46TO57 = 0;
parameter W46TO58 = 0;
parameter W46TO59 = 0;
parameter W46TO60 = 0;
parameter W46TO61 = 0;
parameter W46TO62 = 0;
parameter W46TO63 = 0;
parameter W46TO64 = 0;
parameter W46TO65 = 0;
parameter W46TO66 = 0;
parameter W46TO67 = 0;
parameter W46TO68 = 0;
parameter W46TO69 = 0;
parameter W46TO70 = 0;
parameter W46TO71 = 0;
parameter W46TO72 = 0;
parameter W46TO73 = 0;
parameter W46TO74 = 0;
parameter W46TO75 = 0;
parameter W46TO76 = 0;
parameter W46TO77 = 0;
parameter W46TO78 = 0;
parameter W46TO79 = 0;
parameter W46TO80 = 0;
parameter W46TO81 = 0;
parameter W46TO82 = 0;
parameter W46TO83 = 0;
parameter W46TO84 = 0;
parameter W46TO85 = 0;
parameter W46TO86 = 0;
parameter W46TO87 = 0;
parameter W46TO88 = 0;
parameter W46TO89 = 0;
parameter W46TO90 = 0;
parameter W46TO91 = 0;
parameter W46TO92 = 0;
parameter W46TO93 = 0;
parameter W46TO94 = 0;
parameter W46TO95 = 0;
parameter W46TO96 = 0;
parameter W46TO97 = 0;
parameter W46TO98 = 0;
parameter W46TO99 = 0;
parameter W47TO0 = 0;
parameter W47TO1 = 0;
parameter W47TO2 = 0;
parameter W47TO3 = 0;
parameter W47TO4 = 0;
parameter W47TO5 = 0;
parameter W47TO6 = 0;
parameter W47TO7 = 0;
parameter W47TO8 = 0;
parameter W47TO9 = 0;
parameter W47TO10 = 0;
parameter W47TO11 = 0;
parameter W47TO12 = 0;
parameter W47TO13 = 0;
parameter W47TO14 = 0;
parameter W47TO15 = 0;
parameter W47TO16 = 0;
parameter W47TO17 = 0;
parameter W47TO18 = 0;
parameter W47TO19 = 0;
parameter W47TO20 = 0;
parameter W47TO21 = 0;
parameter W47TO22 = 0;
parameter W47TO23 = 0;
parameter W47TO24 = 0;
parameter W47TO25 = 0;
parameter W47TO26 = 0;
parameter W47TO27 = 0;
parameter W47TO28 = 0;
parameter W47TO29 = 0;
parameter W47TO30 = 0;
parameter W47TO31 = 0;
parameter W47TO32 = 0;
parameter W47TO33 = 0;
parameter W47TO34 = 0;
parameter W47TO35 = 0;
parameter W47TO36 = 0;
parameter W47TO37 = 0;
parameter W47TO38 = 0;
parameter W47TO39 = 0;
parameter W47TO40 = 0;
parameter W47TO41 = 0;
parameter W47TO42 = 0;
parameter W47TO43 = 0;
parameter W47TO44 = 0;
parameter W47TO45 = 0;
parameter W47TO46 = 0;
parameter W47TO47 = 0;
parameter W47TO48 = 0;
parameter W47TO49 = 0;
parameter W47TO50 = 0;
parameter W47TO51 = 0;
parameter W47TO52 = 0;
parameter W47TO53 = 0;
parameter W47TO54 = 0;
parameter W47TO55 = 0;
parameter W47TO56 = 0;
parameter W47TO57 = 0;
parameter W47TO58 = 0;
parameter W47TO59 = 0;
parameter W47TO60 = 0;
parameter W47TO61 = 0;
parameter W47TO62 = 0;
parameter W47TO63 = 0;
parameter W47TO64 = 0;
parameter W47TO65 = 0;
parameter W47TO66 = 0;
parameter W47TO67 = 0;
parameter W47TO68 = 0;
parameter W47TO69 = 0;
parameter W47TO70 = 0;
parameter W47TO71 = 0;
parameter W47TO72 = 0;
parameter W47TO73 = 0;
parameter W47TO74 = 0;
parameter W47TO75 = 0;
parameter W47TO76 = 0;
parameter W47TO77 = 0;
parameter W47TO78 = 0;
parameter W47TO79 = 0;
parameter W47TO80 = 0;
parameter W47TO81 = 0;
parameter W47TO82 = 0;
parameter W47TO83 = 0;
parameter W47TO84 = 0;
parameter W47TO85 = 0;
parameter W47TO86 = 0;
parameter W47TO87 = 0;
parameter W47TO88 = 0;
parameter W47TO89 = 0;
parameter W47TO90 = 0;
parameter W47TO91 = 0;
parameter W47TO92 = 0;
parameter W47TO93 = 0;
parameter W47TO94 = 0;
parameter W47TO95 = 0;
parameter W47TO96 = 0;
parameter W47TO97 = 0;
parameter W47TO98 = 0;
parameter W47TO99 = 0;
parameter W48TO0 = 0;
parameter W48TO1 = 0;
parameter W48TO2 = 0;
parameter W48TO3 = 0;
parameter W48TO4 = 0;
parameter W48TO5 = 0;
parameter W48TO6 = 0;
parameter W48TO7 = 0;
parameter W48TO8 = 0;
parameter W48TO9 = 0;
parameter W48TO10 = 0;
parameter W48TO11 = 0;
parameter W48TO12 = 0;
parameter W48TO13 = 0;
parameter W48TO14 = 0;
parameter W48TO15 = 0;
parameter W48TO16 = 0;
parameter W48TO17 = 0;
parameter W48TO18 = 0;
parameter W48TO19 = 0;
parameter W48TO20 = 0;
parameter W48TO21 = 0;
parameter W48TO22 = 0;
parameter W48TO23 = 0;
parameter W48TO24 = 0;
parameter W48TO25 = 0;
parameter W48TO26 = 0;
parameter W48TO27 = 0;
parameter W48TO28 = 0;
parameter W48TO29 = 0;
parameter W48TO30 = 0;
parameter W48TO31 = 0;
parameter W48TO32 = 0;
parameter W48TO33 = 0;
parameter W48TO34 = 0;
parameter W48TO35 = 0;
parameter W48TO36 = 0;
parameter W48TO37 = 0;
parameter W48TO38 = 0;
parameter W48TO39 = 0;
parameter W48TO40 = 0;
parameter W48TO41 = 0;
parameter W48TO42 = 0;
parameter W48TO43 = 0;
parameter W48TO44 = 0;
parameter W48TO45 = 0;
parameter W48TO46 = 0;
parameter W48TO47 = 0;
parameter W48TO48 = 0;
parameter W48TO49 = 0;
parameter W48TO50 = 0;
parameter W48TO51 = 0;
parameter W48TO52 = 0;
parameter W48TO53 = 0;
parameter W48TO54 = 0;
parameter W48TO55 = 0;
parameter W48TO56 = 0;
parameter W48TO57 = 0;
parameter W48TO58 = 0;
parameter W48TO59 = 0;
parameter W48TO60 = 0;
parameter W48TO61 = 0;
parameter W48TO62 = 0;
parameter W48TO63 = 0;
parameter W48TO64 = 0;
parameter W48TO65 = 0;
parameter W48TO66 = 0;
parameter W48TO67 = 0;
parameter W48TO68 = 0;
parameter W48TO69 = 0;
parameter W48TO70 = 0;
parameter W48TO71 = 0;
parameter W48TO72 = 0;
parameter W48TO73 = 0;
parameter W48TO74 = 0;
parameter W48TO75 = 0;
parameter W48TO76 = 0;
parameter W48TO77 = 0;
parameter W48TO78 = 0;
parameter W48TO79 = 0;
parameter W48TO80 = 0;
parameter W48TO81 = 0;
parameter W48TO82 = 0;
parameter W48TO83 = 0;
parameter W48TO84 = 0;
parameter W48TO85 = 0;
parameter W48TO86 = 0;
parameter W48TO87 = 0;
parameter W48TO88 = 0;
parameter W48TO89 = 0;
parameter W48TO90 = 0;
parameter W48TO91 = 0;
parameter W48TO92 = 0;
parameter W48TO93 = 0;
parameter W48TO94 = 0;
parameter W48TO95 = 0;
parameter W48TO96 = 0;
parameter W48TO97 = 0;
parameter W48TO98 = 0;
parameter W48TO99 = 0;
parameter W49TO0 = 0;
parameter W49TO1 = 0;
parameter W49TO2 = 0;
parameter W49TO3 = 0;
parameter W49TO4 = 0;
parameter W49TO5 = 0;
parameter W49TO6 = 0;
parameter W49TO7 = 0;
parameter W49TO8 = 0;
parameter W49TO9 = 0;
parameter W49TO10 = 0;
parameter W49TO11 = 0;
parameter W49TO12 = 0;
parameter W49TO13 = 0;
parameter W49TO14 = 0;
parameter W49TO15 = 0;
parameter W49TO16 = 0;
parameter W49TO17 = 0;
parameter W49TO18 = 0;
parameter W49TO19 = 0;
parameter W49TO20 = 0;
parameter W49TO21 = 0;
parameter W49TO22 = 0;
parameter W49TO23 = 0;
parameter W49TO24 = 0;
parameter W49TO25 = 0;
parameter W49TO26 = 0;
parameter W49TO27 = 0;
parameter W49TO28 = 0;
parameter W49TO29 = 0;
parameter W49TO30 = 0;
parameter W49TO31 = 0;
parameter W49TO32 = 0;
parameter W49TO33 = 0;
parameter W49TO34 = 0;
parameter W49TO35 = 0;
parameter W49TO36 = 0;
parameter W49TO37 = 0;
parameter W49TO38 = 0;
parameter W49TO39 = 0;
parameter W49TO40 = 0;
parameter W49TO41 = 0;
parameter W49TO42 = 0;
parameter W49TO43 = 0;
parameter W49TO44 = 0;
parameter W49TO45 = 0;
parameter W49TO46 = 0;
parameter W49TO47 = 0;
parameter W49TO48 = 0;
parameter W49TO49 = 0;
parameter W49TO50 = 0;
parameter W49TO51 = 0;
parameter W49TO52 = 0;
parameter W49TO53 = 0;
parameter W49TO54 = 0;
parameter W49TO55 = 0;
parameter W49TO56 = 0;
parameter W49TO57 = 0;
parameter W49TO58 = 0;
parameter W49TO59 = 0;
parameter W49TO60 = 0;
parameter W49TO61 = 0;
parameter W49TO62 = 0;
parameter W49TO63 = 0;
parameter W49TO64 = 0;
parameter W49TO65 = 0;
parameter W49TO66 = 0;
parameter W49TO67 = 0;
parameter W49TO68 = 0;
parameter W49TO69 = 0;
parameter W49TO70 = 0;
parameter W49TO71 = 0;
parameter W49TO72 = 0;
parameter W49TO73 = 0;
parameter W49TO74 = 0;
parameter W49TO75 = 0;
parameter W49TO76 = 0;
parameter W49TO77 = 0;
parameter W49TO78 = 0;
parameter W49TO79 = 0;
parameter W49TO80 = 0;
parameter W49TO81 = 0;
parameter W49TO82 = 0;
parameter W49TO83 = 0;
parameter W49TO84 = 0;
parameter W49TO85 = 0;
parameter W49TO86 = 0;
parameter W49TO87 = 0;
parameter W49TO88 = 0;
parameter W49TO89 = 0;
parameter W49TO90 = 0;
parameter W49TO91 = 0;
parameter W49TO92 = 0;
parameter W49TO93 = 0;
parameter W49TO94 = 0;
parameter W49TO95 = 0;
parameter W49TO96 = 0;
parameter W49TO97 = 0;
parameter W49TO98 = 0;
parameter W49TO99 = 0;
parameter W50TO0 = 0;
parameter W50TO1 = 0;
parameter W50TO2 = 0;
parameter W50TO3 = 0;
parameter W50TO4 = 0;
parameter W50TO5 = 0;
parameter W50TO6 = 0;
parameter W50TO7 = 0;
parameter W50TO8 = 0;
parameter W50TO9 = 0;
parameter W50TO10 = 0;
parameter W50TO11 = 0;
parameter W50TO12 = 0;
parameter W50TO13 = 0;
parameter W50TO14 = 0;
parameter W50TO15 = 0;
parameter W50TO16 = 0;
parameter W50TO17 = 0;
parameter W50TO18 = 0;
parameter W50TO19 = 0;
parameter W50TO20 = 0;
parameter W50TO21 = 0;
parameter W50TO22 = 0;
parameter W50TO23 = 0;
parameter W50TO24 = 0;
parameter W50TO25 = 0;
parameter W50TO26 = 0;
parameter W50TO27 = 0;
parameter W50TO28 = 0;
parameter W50TO29 = 0;
parameter W50TO30 = 0;
parameter W50TO31 = 0;
parameter W50TO32 = 0;
parameter W50TO33 = 0;
parameter W50TO34 = 0;
parameter W50TO35 = 0;
parameter W50TO36 = 0;
parameter W50TO37 = 0;
parameter W50TO38 = 0;
parameter W50TO39 = 0;
parameter W50TO40 = 0;
parameter W50TO41 = 0;
parameter W50TO42 = 0;
parameter W50TO43 = 0;
parameter W50TO44 = 0;
parameter W50TO45 = 0;
parameter W50TO46 = 0;
parameter W50TO47 = 0;
parameter W50TO48 = 0;
parameter W50TO49 = 0;
parameter W50TO50 = 0;
parameter W50TO51 = 0;
parameter W50TO52 = 0;
parameter W50TO53 = 0;
parameter W50TO54 = 0;
parameter W50TO55 = 0;
parameter W50TO56 = 0;
parameter W50TO57 = 0;
parameter W50TO58 = 0;
parameter W50TO59 = 0;
parameter W50TO60 = 0;
parameter W50TO61 = 0;
parameter W50TO62 = 0;
parameter W50TO63 = 0;
parameter W50TO64 = 0;
parameter W50TO65 = 0;
parameter W50TO66 = 0;
parameter W50TO67 = 0;
parameter W50TO68 = 0;
parameter W50TO69 = 0;
parameter W50TO70 = 0;
parameter W50TO71 = 0;
parameter W50TO72 = 0;
parameter W50TO73 = 0;
parameter W50TO74 = 0;
parameter W50TO75 = 0;
parameter W50TO76 = 0;
parameter W50TO77 = 0;
parameter W50TO78 = 0;
parameter W50TO79 = 0;
parameter W50TO80 = 0;
parameter W50TO81 = 0;
parameter W50TO82 = 0;
parameter W50TO83 = 0;
parameter W50TO84 = 0;
parameter W50TO85 = 0;
parameter W50TO86 = 0;
parameter W50TO87 = 0;
parameter W50TO88 = 0;
parameter W50TO89 = 0;
parameter W50TO90 = 0;
parameter W50TO91 = 0;
parameter W50TO92 = 0;
parameter W50TO93 = 0;
parameter W50TO94 = 0;
parameter W50TO95 = 0;
parameter W50TO96 = 0;
parameter W50TO97 = 0;
parameter W50TO98 = 0;
parameter W50TO99 = 0;
parameter W51TO0 = 0;
parameter W51TO1 = 0;
parameter W51TO2 = 0;
parameter W51TO3 = 0;
parameter W51TO4 = 0;
parameter W51TO5 = 0;
parameter W51TO6 = 0;
parameter W51TO7 = 0;
parameter W51TO8 = 0;
parameter W51TO9 = 0;
parameter W51TO10 = 0;
parameter W51TO11 = 0;
parameter W51TO12 = 0;
parameter W51TO13 = 0;
parameter W51TO14 = 0;
parameter W51TO15 = 0;
parameter W51TO16 = 0;
parameter W51TO17 = 0;
parameter W51TO18 = 0;
parameter W51TO19 = 0;
parameter W51TO20 = 0;
parameter W51TO21 = 0;
parameter W51TO22 = 0;
parameter W51TO23 = 0;
parameter W51TO24 = 0;
parameter W51TO25 = 0;
parameter W51TO26 = 0;
parameter W51TO27 = 0;
parameter W51TO28 = 0;
parameter W51TO29 = 0;
parameter W51TO30 = 0;
parameter W51TO31 = 0;
parameter W51TO32 = 0;
parameter W51TO33 = 0;
parameter W51TO34 = 0;
parameter W51TO35 = 0;
parameter W51TO36 = 0;
parameter W51TO37 = 0;
parameter W51TO38 = 0;
parameter W51TO39 = 0;
parameter W51TO40 = 0;
parameter W51TO41 = 0;
parameter W51TO42 = 0;
parameter W51TO43 = 0;
parameter W51TO44 = 0;
parameter W51TO45 = 0;
parameter W51TO46 = 0;
parameter W51TO47 = 0;
parameter W51TO48 = 0;
parameter W51TO49 = 0;
parameter W51TO50 = 0;
parameter W51TO51 = 0;
parameter W51TO52 = 0;
parameter W51TO53 = 0;
parameter W51TO54 = 0;
parameter W51TO55 = 0;
parameter W51TO56 = 0;
parameter W51TO57 = 0;
parameter W51TO58 = 0;
parameter W51TO59 = 0;
parameter W51TO60 = 0;
parameter W51TO61 = 0;
parameter W51TO62 = 0;
parameter W51TO63 = 0;
parameter W51TO64 = 0;
parameter W51TO65 = 0;
parameter W51TO66 = 0;
parameter W51TO67 = 0;
parameter W51TO68 = 0;
parameter W51TO69 = 0;
parameter W51TO70 = 0;
parameter W51TO71 = 0;
parameter W51TO72 = 0;
parameter W51TO73 = 0;
parameter W51TO74 = 0;
parameter W51TO75 = 0;
parameter W51TO76 = 0;
parameter W51TO77 = 0;
parameter W51TO78 = 0;
parameter W51TO79 = 0;
parameter W51TO80 = 0;
parameter W51TO81 = 0;
parameter W51TO82 = 0;
parameter W51TO83 = 0;
parameter W51TO84 = 0;
parameter W51TO85 = 0;
parameter W51TO86 = 0;
parameter W51TO87 = 0;
parameter W51TO88 = 0;
parameter W51TO89 = 0;
parameter W51TO90 = 0;
parameter W51TO91 = 0;
parameter W51TO92 = 0;
parameter W51TO93 = 0;
parameter W51TO94 = 0;
parameter W51TO95 = 0;
parameter W51TO96 = 0;
parameter W51TO97 = 0;
parameter W51TO98 = 0;
parameter W51TO99 = 0;
parameter W52TO0 = 0;
parameter W52TO1 = 0;
parameter W52TO2 = 0;
parameter W52TO3 = 0;
parameter W52TO4 = 0;
parameter W52TO5 = 0;
parameter W52TO6 = 0;
parameter W52TO7 = 0;
parameter W52TO8 = 0;
parameter W52TO9 = 0;
parameter W52TO10 = 0;
parameter W52TO11 = 0;
parameter W52TO12 = 0;
parameter W52TO13 = 0;
parameter W52TO14 = 0;
parameter W52TO15 = 0;
parameter W52TO16 = 0;
parameter W52TO17 = 0;
parameter W52TO18 = 0;
parameter W52TO19 = 0;
parameter W52TO20 = 0;
parameter W52TO21 = 0;
parameter W52TO22 = 0;
parameter W52TO23 = 0;
parameter W52TO24 = 0;
parameter W52TO25 = 0;
parameter W52TO26 = 0;
parameter W52TO27 = 0;
parameter W52TO28 = 0;
parameter W52TO29 = 0;
parameter W52TO30 = 0;
parameter W52TO31 = 0;
parameter W52TO32 = 0;
parameter W52TO33 = 0;
parameter W52TO34 = 0;
parameter W52TO35 = 0;
parameter W52TO36 = 0;
parameter W52TO37 = 0;
parameter W52TO38 = 0;
parameter W52TO39 = 0;
parameter W52TO40 = 0;
parameter W52TO41 = 0;
parameter W52TO42 = 0;
parameter W52TO43 = 0;
parameter W52TO44 = 0;
parameter W52TO45 = 0;
parameter W52TO46 = 0;
parameter W52TO47 = 0;
parameter W52TO48 = 0;
parameter W52TO49 = 0;
parameter W52TO50 = 0;
parameter W52TO51 = 0;
parameter W52TO52 = 0;
parameter W52TO53 = 0;
parameter W52TO54 = 0;
parameter W52TO55 = 0;
parameter W52TO56 = 0;
parameter W52TO57 = 0;
parameter W52TO58 = 0;
parameter W52TO59 = 0;
parameter W52TO60 = 0;
parameter W52TO61 = 0;
parameter W52TO62 = 0;
parameter W52TO63 = 0;
parameter W52TO64 = 0;
parameter W52TO65 = 0;
parameter W52TO66 = 0;
parameter W52TO67 = 0;
parameter W52TO68 = 0;
parameter W52TO69 = 0;
parameter W52TO70 = 0;
parameter W52TO71 = 0;
parameter W52TO72 = 0;
parameter W52TO73 = 0;
parameter W52TO74 = 0;
parameter W52TO75 = 0;
parameter W52TO76 = 0;
parameter W52TO77 = 0;
parameter W52TO78 = 0;
parameter W52TO79 = 0;
parameter W52TO80 = 0;
parameter W52TO81 = 0;
parameter W52TO82 = 0;
parameter W52TO83 = 0;
parameter W52TO84 = 0;
parameter W52TO85 = 0;
parameter W52TO86 = 0;
parameter W52TO87 = 0;
parameter W52TO88 = 0;
parameter W52TO89 = 0;
parameter W52TO90 = 0;
parameter W52TO91 = 0;
parameter W52TO92 = 0;
parameter W52TO93 = 0;
parameter W52TO94 = 0;
parameter W52TO95 = 0;
parameter W52TO96 = 0;
parameter W52TO97 = 0;
parameter W52TO98 = 0;
parameter W52TO99 = 0;
parameter W53TO0 = 0;
parameter W53TO1 = 0;
parameter W53TO2 = 0;
parameter W53TO3 = 0;
parameter W53TO4 = 0;
parameter W53TO5 = 0;
parameter W53TO6 = 0;
parameter W53TO7 = 0;
parameter W53TO8 = 0;
parameter W53TO9 = 0;
parameter W53TO10 = 0;
parameter W53TO11 = 0;
parameter W53TO12 = 0;
parameter W53TO13 = 0;
parameter W53TO14 = 0;
parameter W53TO15 = 0;
parameter W53TO16 = 0;
parameter W53TO17 = 0;
parameter W53TO18 = 0;
parameter W53TO19 = 0;
parameter W53TO20 = 0;
parameter W53TO21 = 0;
parameter W53TO22 = 0;
parameter W53TO23 = 0;
parameter W53TO24 = 0;
parameter W53TO25 = 0;
parameter W53TO26 = 0;
parameter W53TO27 = 0;
parameter W53TO28 = 0;
parameter W53TO29 = 0;
parameter W53TO30 = 0;
parameter W53TO31 = 0;
parameter W53TO32 = 0;
parameter W53TO33 = 0;
parameter W53TO34 = 0;
parameter W53TO35 = 0;
parameter W53TO36 = 0;
parameter W53TO37 = 0;
parameter W53TO38 = 0;
parameter W53TO39 = 0;
parameter W53TO40 = 0;
parameter W53TO41 = 0;
parameter W53TO42 = 0;
parameter W53TO43 = 0;
parameter W53TO44 = 0;
parameter W53TO45 = 0;
parameter W53TO46 = 0;
parameter W53TO47 = 0;
parameter W53TO48 = 0;
parameter W53TO49 = 0;
parameter W53TO50 = 0;
parameter W53TO51 = 0;
parameter W53TO52 = 0;
parameter W53TO53 = 0;
parameter W53TO54 = 0;
parameter W53TO55 = 0;
parameter W53TO56 = 0;
parameter W53TO57 = 0;
parameter W53TO58 = 0;
parameter W53TO59 = 0;
parameter W53TO60 = 0;
parameter W53TO61 = 0;
parameter W53TO62 = 0;
parameter W53TO63 = 0;
parameter W53TO64 = 0;
parameter W53TO65 = 0;
parameter W53TO66 = 0;
parameter W53TO67 = 0;
parameter W53TO68 = 0;
parameter W53TO69 = 0;
parameter W53TO70 = 0;
parameter W53TO71 = 0;
parameter W53TO72 = 0;
parameter W53TO73 = 0;
parameter W53TO74 = 0;
parameter W53TO75 = 0;
parameter W53TO76 = 0;
parameter W53TO77 = 0;
parameter W53TO78 = 0;
parameter W53TO79 = 0;
parameter W53TO80 = 0;
parameter W53TO81 = 0;
parameter W53TO82 = 0;
parameter W53TO83 = 0;
parameter W53TO84 = 0;
parameter W53TO85 = 0;
parameter W53TO86 = 0;
parameter W53TO87 = 0;
parameter W53TO88 = 0;
parameter W53TO89 = 0;
parameter W53TO90 = 0;
parameter W53TO91 = 0;
parameter W53TO92 = 0;
parameter W53TO93 = 0;
parameter W53TO94 = 0;
parameter W53TO95 = 0;
parameter W53TO96 = 0;
parameter W53TO97 = 0;
parameter W53TO98 = 0;
parameter W53TO99 = 0;
parameter W54TO0 = 0;
parameter W54TO1 = 0;
parameter W54TO2 = 0;
parameter W54TO3 = 0;
parameter W54TO4 = 0;
parameter W54TO5 = 0;
parameter W54TO6 = 0;
parameter W54TO7 = 0;
parameter W54TO8 = 0;
parameter W54TO9 = 0;
parameter W54TO10 = 0;
parameter W54TO11 = 0;
parameter W54TO12 = 0;
parameter W54TO13 = 0;
parameter W54TO14 = 0;
parameter W54TO15 = 0;
parameter W54TO16 = 0;
parameter W54TO17 = 0;
parameter W54TO18 = 0;
parameter W54TO19 = 0;
parameter W54TO20 = 0;
parameter W54TO21 = 0;
parameter W54TO22 = 0;
parameter W54TO23 = 0;
parameter W54TO24 = 0;
parameter W54TO25 = 0;
parameter W54TO26 = 0;
parameter W54TO27 = 0;
parameter W54TO28 = 0;
parameter W54TO29 = 0;
parameter W54TO30 = 0;
parameter W54TO31 = 0;
parameter W54TO32 = 0;
parameter W54TO33 = 0;
parameter W54TO34 = 0;
parameter W54TO35 = 0;
parameter W54TO36 = 0;
parameter W54TO37 = 0;
parameter W54TO38 = 0;
parameter W54TO39 = 0;
parameter W54TO40 = 0;
parameter W54TO41 = 0;
parameter W54TO42 = 0;
parameter W54TO43 = 0;
parameter W54TO44 = 0;
parameter W54TO45 = 0;
parameter W54TO46 = 0;
parameter W54TO47 = 0;
parameter W54TO48 = 0;
parameter W54TO49 = 0;
parameter W54TO50 = 0;
parameter W54TO51 = 0;
parameter W54TO52 = 0;
parameter W54TO53 = 0;
parameter W54TO54 = 0;
parameter W54TO55 = 0;
parameter W54TO56 = 0;
parameter W54TO57 = 0;
parameter W54TO58 = 0;
parameter W54TO59 = 0;
parameter W54TO60 = 0;
parameter W54TO61 = 0;
parameter W54TO62 = 0;
parameter W54TO63 = 0;
parameter W54TO64 = 0;
parameter W54TO65 = 0;
parameter W54TO66 = 0;
parameter W54TO67 = 0;
parameter W54TO68 = 0;
parameter W54TO69 = 0;
parameter W54TO70 = 0;
parameter W54TO71 = 0;
parameter W54TO72 = 0;
parameter W54TO73 = 0;
parameter W54TO74 = 0;
parameter W54TO75 = 0;
parameter W54TO76 = 0;
parameter W54TO77 = 0;
parameter W54TO78 = 0;
parameter W54TO79 = 0;
parameter W54TO80 = 0;
parameter W54TO81 = 0;
parameter W54TO82 = 0;
parameter W54TO83 = 0;
parameter W54TO84 = 0;
parameter W54TO85 = 0;
parameter W54TO86 = 0;
parameter W54TO87 = 0;
parameter W54TO88 = 0;
parameter W54TO89 = 0;
parameter W54TO90 = 0;
parameter W54TO91 = 0;
parameter W54TO92 = 0;
parameter W54TO93 = 0;
parameter W54TO94 = 0;
parameter W54TO95 = 0;
parameter W54TO96 = 0;
parameter W54TO97 = 0;
parameter W54TO98 = 0;
parameter W54TO99 = 0;
parameter W55TO0 = 0;
parameter W55TO1 = 0;
parameter W55TO2 = 0;
parameter W55TO3 = 0;
parameter W55TO4 = 0;
parameter W55TO5 = 0;
parameter W55TO6 = 0;
parameter W55TO7 = 0;
parameter W55TO8 = 0;
parameter W55TO9 = 0;
parameter W55TO10 = 0;
parameter W55TO11 = 0;
parameter W55TO12 = 0;
parameter W55TO13 = 0;
parameter W55TO14 = 0;
parameter W55TO15 = 0;
parameter W55TO16 = 0;
parameter W55TO17 = 0;
parameter W55TO18 = 0;
parameter W55TO19 = 0;
parameter W55TO20 = 0;
parameter W55TO21 = 0;
parameter W55TO22 = 0;
parameter W55TO23 = 0;
parameter W55TO24 = 0;
parameter W55TO25 = 0;
parameter W55TO26 = 0;
parameter W55TO27 = 0;
parameter W55TO28 = 0;
parameter W55TO29 = 0;
parameter W55TO30 = 0;
parameter W55TO31 = 0;
parameter W55TO32 = 0;
parameter W55TO33 = 0;
parameter W55TO34 = 0;
parameter W55TO35 = 0;
parameter W55TO36 = 0;
parameter W55TO37 = 0;
parameter W55TO38 = 0;
parameter W55TO39 = 0;
parameter W55TO40 = 0;
parameter W55TO41 = 0;
parameter W55TO42 = 0;
parameter W55TO43 = 0;
parameter W55TO44 = 0;
parameter W55TO45 = 0;
parameter W55TO46 = 0;
parameter W55TO47 = 0;
parameter W55TO48 = 0;
parameter W55TO49 = 0;
parameter W55TO50 = 0;
parameter W55TO51 = 0;
parameter W55TO52 = 0;
parameter W55TO53 = 0;
parameter W55TO54 = 0;
parameter W55TO55 = 0;
parameter W55TO56 = 0;
parameter W55TO57 = 0;
parameter W55TO58 = 0;
parameter W55TO59 = 0;
parameter W55TO60 = 0;
parameter W55TO61 = 0;
parameter W55TO62 = 0;
parameter W55TO63 = 0;
parameter W55TO64 = 0;
parameter W55TO65 = 0;
parameter W55TO66 = 0;
parameter W55TO67 = 0;
parameter W55TO68 = 0;
parameter W55TO69 = 0;
parameter W55TO70 = 0;
parameter W55TO71 = 0;
parameter W55TO72 = 0;
parameter W55TO73 = 0;
parameter W55TO74 = 0;
parameter W55TO75 = 0;
parameter W55TO76 = 0;
parameter W55TO77 = 0;
parameter W55TO78 = 0;
parameter W55TO79 = 0;
parameter W55TO80 = 0;
parameter W55TO81 = 0;
parameter W55TO82 = 0;
parameter W55TO83 = 0;
parameter W55TO84 = 0;
parameter W55TO85 = 0;
parameter W55TO86 = 0;
parameter W55TO87 = 0;
parameter W55TO88 = 0;
parameter W55TO89 = 0;
parameter W55TO90 = 0;
parameter W55TO91 = 0;
parameter W55TO92 = 0;
parameter W55TO93 = 0;
parameter W55TO94 = 0;
parameter W55TO95 = 0;
parameter W55TO96 = 0;
parameter W55TO97 = 0;
parameter W55TO98 = 0;
parameter W55TO99 = 0;
parameter W56TO0 = 0;
parameter W56TO1 = 0;
parameter W56TO2 = 0;
parameter W56TO3 = 0;
parameter W56TO4 = 0;
parameter W56TO5 = 0;
parameter W56TO6 = 0;
parameter W56TO7 = 0;
parameter W56TO8 = 0;
parameter W56TO9 = 0;
parameter W56TO10 = 0;
parameter W56TO11 = 0;
parameter W56TO12 = 0;
parameter W56TO13 = 0;
parameter W56TO14 = 0;
parameter W56TO15 = 0;
parameter W56TO16 = 0;
parameter W56TO17 = 0;
parameter W56TO18 = 0;
parameter W56TO19 = 0;
parameter W56TO20 = 0;
parameter W56TO21 = 0;
parameter W56TO22 = 0;
parameter W56TO23 = 0;
parameter W56TO24 = 0;
parameter W56TO25 = 0;
parameter W56TO26 = 0;
parameter W56TO27 = 0;
parameter W56TO28 = 0;
parameter W56TO29 = 0;
parameter W56TO30 = 0;
parameter W56TO31 = 0;
parameter W56TO32 = 0;
parameter W56TO33 = 0;
parameter W56TO34 = 0;
parameter W56TO35 = 0;
parameter W56TO36 = 0;
parameter W56TO37 = 0;
parameter W56TO38 = 0;
parameter W56TO39 = 0;
parameter W56TO40 = 0;
parameter W56TO41 = 0;
parameter W56TO42 = 0;
parameter W56TO43 = 0;
parameter W56TO44 = 0;
parameter W56TO45 = 0;
parameter W56TO46 = 0;
parameter W56TO47 = 0;
parameter W56TO48 = 0;
parameter W56TO49 = 0;
parameter W56TO50 = 0;
parameter W56TO51 = 0;
parameter W56TO52 = 0;
parameter W56TO53 = 0;
parameter W56TO54 = 0;
parameter W56TO55 = 0;
parameter W56TO56 = 0;
parameter W56TO57 = 0;
parameter W56TO58 = 0;
parameter W56TO59 = 0;
parameter W56TO60 = 0;
parameter W56TO61 = 0;
parameter W56TO62 = 0;
parameter W56TO63 = 0;
parameter W56TO64 = 0;
parameter W56TO65 = 0;
parameter W56TO66 = 0;
parameter W56TO67 = 0;
parameter W56TO68 = 0;
parameter W56TO69 = 0;
parameter W56TO70 = 0;
parameter W56TO71 = 0;
parameter W56TO72 = 0;
parameter W56TO73 = 0;
parameter W56TO74 = 0;
parameter W56TO75 = 0;
parameter W56TO76 = 0;
parameter W56TO77 = 0;
parameter W56TO78 = 0;
parameter W56TO79 = 0;
parameter W56TO80 = 0;
parameter W56TO81 = 0;
parameter W56TO82 = 0;
parameter W56TO83 = 0;
parameter W56TO84 = 0;
parameter W56TO85 = 0;
parameter W56TO86 = 0;
parameter W56TO87 = 0;
parameter W56TO88 = 0;
parameter W56TO89 = 0;
parameter W56TO90 = 0;
parameter W56TO91 = 0;
parameter W56TO92 = 0;
parameter W56TO93 = 0;
parameter W56TO94 = 0;
parameter W56TO95 = 0;
parameter W56TO96 = 0;
parameter W56TO97 = 0;
parameter W56TO98 = 0;
parameter W56TO99 = 0;
parameter W57TO0 = 0;
parameter W57TO1 = 0;
parameter W57TO2 = 0;
parameter W57TO3 = 0;
parameter W57TO4 = 0;
parameter W57TO5 = 0;
parameter W57TO6 = 0;
parameter W57TO7 = 0;
parameter W57TO8 = 0;
parameter W57TO9 = 0;
parameter W57TO10 = 0;
parameter W57TO11 = 0;
parameter W57TO12 = 0;
parameter W57TO13 = 0;
parameter W57TO14 = 0;
parameter W57TO15 = 0;
parameter W57TO16 = 0;
parameter W57TO17 = 0;
parameter W57TO18 = 0;
parameter W57TO19 = 0;
parameter W57TO20 = 0;
parameter W57TO21 = 0;
parameter W57TO22 = 0;
parameter W57TO23 = 0;
parameter W57TO24 = 0;
parameter W57TO25 = 0;
parameter W57TO26 = 0;
parameter W57TO27 = 0;
parameter W57TO28 = 0;
parameter W57TO29 = 0;
parameter W57TO30 = 0;
parameter W57TO31 = 0;
parameter W57TO32 = 0;
parameter W57TO33 = 0;
parameter W57TO34 = 0;
parameter W57TO35 = 0;
parameter W57TO36 = 0;
parameter W57TO37 = 0;
parameter W57TO38 = 0;
parameter W57TO39 = 0;
parameter W57TO40 = 0;
parameter W57TO41 = 0;
parameter W57TO42 = 0;
parameter W57TO43 = 0;
parameter W57TO44 = 0;
parameter W57TO45 = 0;
parameter W57TO46 = 0;
parameter W57TO47 = 0;
parameter W57TO48 = 0;
parameter W57TO49 = 0;
parameter W57TO50 = 0;
parameter W57TO51 = 0;
parameter W57TO52 = 0;
parameter W57TO53 = 0;
parameter W57TO54 = 0;
parameter W57TO55 = 0;
parameter W57TO56 = 0;
parameter W57TO57 = 0;
parameter W57TO58 = 0;
parameter W57TO59 = 0;
parameter W57TO60 = 0;
parameter W57TO61 = 0;
parameter W57TO62 = 0;
parameter W57TO63 = 0;
parameter W57TO64 = 0;
parameter W57TO65 = 0;
parameter W57TO66 = 0;
parameter W57TO67 = 0;
parameter W57TO68 = 0;
parameter W57TO69 = 0;
parameter W57TO70 = 0;
parameter W57TO71 = 0;
parameter W57TO72 = 0;
parameter W57TO73 = 0;
parameter W57TO74 = 0;
parameter W57TO75 = 0;
parameter W57TO76 = 0;
parameter W57TO77 = 0;
parameter W57TO78 = 0;
parameter W57TO79 = 0;
parameter W57TO80 = 0;
parameter W57TO81 = 0;
parameter W57TO82 = 0;
parameter W57TO83 = 0;
parameter W57TO84 = 0;
parameter W57TO85 = 0;
parameter W57TO86 = 0;
parameter W57TO87 = 0;
parameter W57TO88 = 0;
parameter W57TO89 = 0;
parameter W57TO90 = 0;
parameter W57TO91 = 0;
parameter W57TO92 = 0;
parameter W57TO93 = 0;
parameter W57TO94 = 0;
parameter W57TO95 = 0;
parameter W57TO96 = 0;
parameter W57TO97 = 0;
parameter W57TO98 = 0;
parameter W57TO99 = 0;
parameter W58TO0 = 0;
parameter W58TO1 = 0;
parameter W58TO2 = 0;
parameter W58TO3 = 0;
parameter W58TO4 = 0;
parameter W58TO5 = 0;
parameter W58TO6 = 0;
parameter W58TO7 = 0;
parameter W58TO8 = 0;
parameter W58TO9 = 0;
parameter W58TO10 = 0;
parameter W58TO11 = 0;
parameter W58TO12 = 0;
parameter W58TO13 = 0;
parameter W58TO14 = 0;
parameter W58TO15 = 0;
parameter W58TO16 = 0;
parameter W58TO17 = 0;
parameter W58TO18 = 0;
parameter W58TO19 = 0;
parameter W58TO20 = 0;
parameter W58TO21 = 0;
parameter W58TO22 = 0;
parameter W58TO23 = 0;
parameter W58TO24 = 0;
parameter W58TO25 = 0;
parameter W58TO26 = 0;
parameter W58TO27 = 0;
parameter W58TO28 = 0;
parameter W58TO29 = 0;
parameter W58TO30 = 0;
parameter W58TO31 = 0;
parameter W58TO32 = 0;
parameter W58TO33 = 0;
parameter W58TO34 = 0;
parameter W58TO35 = 0;
parameter W58TO36 = 0;
parameter W58TO37 = 0;
parameter W58TO38 = 0;
parameter W58TO39 = 0;
parameter W58TO40 = 0;
parameter W58TO41 = 0;
parameter W58TO42 = 0;
parameter W58TO43 = 0;
parameter W58TO44 = 0;
parameter W58TO45 = 0;
parameter W58TO46 = 0;
parameter W58TO47 = 0;
parameter W58TO48 = 0;
parameter W58TO49 = 0;
parameter W58TO50 = 0;
parameter W58TO51 = 0;
parameter W58TO52 = 0;
parameter W58TO53 = 0;
parameter W58TO54 = 0;
parameter W58TO55 = 0;
parameter W58TO56 = 0;
parameter W58TO57 = 0;
parameter W58TO58 = 0;
parameter W58TO59 = 0;
parameter W58TO60 = 0;
parameter W58TO61 = 0;
parameter W58TO62 = 0;
parameter W58TO63 = 0;
parameter W58TO64 = 0;
parameter W58TO65 = 0;
parameter W58TO66 = 0;
parameter W58TO67 = 0;
parameter W58TO68 = 0;
parameter W58TO69 = 0;
parameter W58TO70 = 0;
parameter W58TO71 = 0;
parameter W58TO72 = 0;
parameter W58TO73 = 0;
parameter W58TO74 = 0;
parameter W58TO75 = 0;
parameter W58TO76 = 0;
parameter W58TO77 = 0;
parameter W58TO78 = 0;
parameter W58TO79 = 0;
parameter W58TO80 = 0;
parameter W58TO81 = 0;
parameter W58TO82 = 0;
parameter W58TO83 = 0;
parameter W58TO84 = 0;
parameter W58TO85 = 0;
parameter W58TO86 = 0;
parameter W58TO87 = 0;
parameter W58TO88 = 0;
parameter W58TO89 = 0;
parameter W58TO90 = 0;
parameter W58TO91 = 0;
parameter W58TO92 = 0;
parameter W58TO93 = 0;
parameter W58TO94 = 0;
parameter W58TO95 = 0;
parameter W58TO96 = 0;
parameter W58TO97 = 0;
parameter W58TO98 = 0;
parameter W58TO99 = 0;
parameter W59TO0 = 0;
parameter W59TO1 = 0;
parameter W59TO2 = 0;
parameter W59TO3 = 0;
parameter W59TO4 = 0;
parameter W59TO5 = 0;
parameter W59TO6 = 0;
parameter W59TO7 = 0;
parameter W59TO8 = 0;
parameter W59TO9 = 0;
parameter W59TO10 = 0;
parameter W59TO11 = 0;
parameter W59TO12 = 0;
parameter W59TO13 = 0;
parameter W59TO14 = 0;
parameter W59TO15 = 0;
parameter W59TO16 = 0;
parameter W59TO17 = 0;
parameter W59TO18 = 0;
parameter W59TO19 = 0;
parameter W59TO20 = 0;
parameter W59TO21 = 0;
parameter W59TO22 = 0;
parameter W59TO23 = 0;
parameter W59TO24 = 0;
parameter W59TO25 = 0;
parameter W59TO26 = 0;
parameter W59TO27 = 0;
parameter W59TO28 = 0;
parameter W59TO29 = 0;
parameter W59TO30 = 0;
parameter W59TO31 = 0;
parameter W59TO32 = 0;
parameter W59TO33 = 0;
parameter W59TO34 = 0;
parameter W59TO35 = 0;
parameter W59TO36 = 0;
parameter W59TO37 = 0;
parameter W59TO38 = 0;
parameter W59TO39 = 0;
parameter W59TO40 = 0;
parameter W59TO41 = 0;
parameter W59TO42 = 0;
parameter W59TO43 = 0;
parameter W59TO44 = 0;
parameter W59TO45 = 0;
parameter W59TO46 = 0;
parameter W59TO47 = 0;
parameter W59TO48 = 0;
parameter W59TO49 = 0;
parameter W59TO50 = 0;
parameter W59TO51 = 0;
parameter W59TO52 = 0;
parameter W59TO53 = 0;
parameter W59TO54 = 0;
parameter W59TO55 = 0;
parameter W59TO56 = 0;
parameter W59TO57 = 0;
parameter W59TO58 = 0;
parameter W59TO59 = 0;
parameter W59TO60 = 0;
parameter W59TO61 = 0;
parameter W59TO62 = 0;
parameter W59TO63 = 0;
parameter W59TO64 = 0;
parameter W59TO65 = 0;
parameter W59TO66 = 0;
parameter W59TO67 = 0;
parameter W59TO68 = 0;
parameter W59TO69 = 0;
parameter W59TO70 = 0;
parameter W59TO71 = 0;
parameter W59TO72 = 0;
parameter W59TO73 = 0;
parameter W59TO74 = 0;
parameter W59TO75 = 0;
parameter W59TO76 = 0;
parameter W59TO77 = 0;
parameter W59TO78 = 0;
parameter W59TO79 = 0;
parameter W59TO80 = 0;
parameter W59TO81 = 0;
parameter W59TO82 = 0;
parameter W59TO83 = 0;
parameter W59TO84 = 0;
parameter W59TO85 = 0;
parameter W59TO86 = 0;
parameter W59TO87 = 0;
parameter W59TO88 = 0;
parameter W59TO89 = 0;
parameter W59TO90 = 0;
parameter W59TO91 = 0;
parameter W59TO92 = 0;
parameter W59TO93 = 0;
parameter W59TO94 = 0;
parameter W59TO95 = 0;
parameter W59TO96 = 0;
parameter W59TO97 = 0;
parameter W59TO98 = 0;
parameter W59TO99 = 0;
parameter W60TO0 = 0;
parameter W60TO1 = 0;
parameter W60TO2 = 0;
parameter W60TO3 = 0;
parameter W60TO4 = 0;
parameter W60TO5 = 0;
parameter W60TO6 = 0;
parameter W60TO7 = 0;
parameter W60TO8 = 0;
parameter W60TO9 = 0;
parameter W60TO10 = 0;
parameter W60TO11 = 0;
parameter W60TO12 = 0;
parameter W60TO13 = 0;
parameter W60TO14 = 0;
parameter W60TO15 = 0;
parameter W60TO16 = 0;
parameter W60TO17 = 0;
parameter W60TO18 = 0;
parameter W60TO19 = 0;
parameter W60TO20 = 0;
parameter W60TO21 = 0;
parameter W60TO22 = 0;
parameter W60TO23 = 0;
parameter W60TO24 = 0;
parameter W60TO25 = 0;
parameter W60TO26 = 0;
parameter W60TO27 = 0;
parameter W60TO28 = 0;
parameter W60TO29 = 0;
parameter W60TO30 = 0;
parameter W60TO31 = 0;
parameter W60TO32 = 0;
parameter W60TO33 = 0;
parameter W60TO34 = 0;
parameter W60TO35 = 0;
parameter W60TO36 = 0;
parameter W60TO37 = 0;
parameter W60TO38 = 0;
parameter W60TO39 = 0;
parameter W60TO40 = 0;
parameter W60TO41 = 0;
parameter W60TO42 = 0;
parameter W60TO43 = 0;
parameter W60TO44 = 0;
parameter W60TO45 = 0;
parameter W60TO46 = 0;
parameter W60TO47 = 0;
parameter W60TO48 = 0;
parameter W60TO49 = 0;
parameter W60TO50 = 0;
parameter W60TO51 = 0;
parameter W60TO52 = 0;
parameter W60TO53 = 0;
parameter W60TO54 = 0;
parameter W60TO55 = 0;
parameter W60TO56 = 0;
parameter W60TO57 = 0;
parameter W60TO58 = 0;
parameter W60TO59 = 0;
parameter W60TO60 = 0;
parameter W60TO61 = 0;
parameter W60TO62 = 0;
parameter W60TO63 = 0;
parameter W60TO64 = 0;
parameter W60TO65 = 0;
parameter W60TO66 = 0;
parameter W60TO67 = 0;
parameter W60TO68 = 0;
parameter W60TO69 = 0;
parameter W60TO70 = 0;
parameter W60TO71 = 0;
parameter W60TO72 = 0;
parameter W60TO73 = 0;
parameter W60TO74 = 0;
parameter W60TO75 = 0;
parameter W60TO76 = 0;
parameter W60TO77 = 0;
parameter W60TO78 = 0;
parameter W60TO79 = 0;
parameter W60TO80 = 0;
parameter W60TO81 = 0;
parameter W60TO82 = 0;
parameter W60TO83 = 0;
parameter W60TO84 = 0;
parameter W60TO85 = 0;
parameter W60TO86 = 0;
parameter W60TO87 = 0;
parameter W60TO88 = 0;
parameter W60TO89 = 0;
parameter W60TO90 = 0;
parameter W60TO91 = 0;
parameter W60TO92 = 0;
parameter W60TO93 = 0;
parameter W60TO94 = 0;
parameter W60TO95 = 0;
parameter W60TO96 = 0;
parameter W60TO97 = 0;
parameter W60TO98 = 0;
parameter W60TO99 = 0;
parameter W61TO0 = 0;
parameter W61TO1 = 0;
parameter W61TO2 = 0;
parameter W61TO3 = 0;
parameter W61TO4 = 0;
parameter W61TO5 = 0;
parameter W61TO6 = 0;
parameter W61TO7 = 0;
parameter W61TO8 = 0;
parameter W61TO9 = 0;
parameter W61TO10 = 0;
parameter W61TO11 = 0;
parameter W61TO12 = 0;
parameter W61TO13 = 0;
parameter W61TO14 = 0;
parameter W61TO15 = 0;
parameter W61TO16 = 0;
parameter W61TO17 = 0;
parameter W61TO18 = 0;
parameter W61TO19 = 0;
parameter W61TO20 = 0;
parameter W61TO21 = 0;
parameter W61TO22 = 0;
parameter W61TO23 = 0;
parameter W61TO24 = 0;
parameter W61TO25 = 0;
parameter W61TO26 = 0;
parameter W61TO27 = 0;
parameter W61TO28 = 0;
parameter W61TO29 = 0;
parameter W61TO30 = 0;
parameter W61TO31 = 0;
parameter W61TO32 = 0;
parameter W61TO33 = 0;
parameter W61TO34 = 0;
parameter W61TO35 = 0;
parameter W61TO36 = 0;
parameter W61TO37 = 0;
parameter W61TO38 = 0;
parameter W61TO39 = 0;
parameter W61TO40 = 0;
parameter W61TO41 = 0;
parameter W61TO42 = 0;
parameter W61TO43 = 0;
parameter W61TO44 = 0;
parameter W61TO45 = 0;
parameter W61TO46 = 0;
parameter W61TO47 = 0;
parameter W61TO48 = 0;
parameter W61TO49 = 0;
parameter W61TO50 = 0;
parameter W61TO51 = 0;
parameter W61TO52 = 0;
parameter W61TO53 = 0;
parameter W61TO54 = 0;
parameter W61TO55 = 0;
parameter W61TO56 = 0;
parameter W61TO57 = 0;
parameter W61TO58 = 0;
parameter W61TO59 = 0;
parameter W61TO60 = 0;
parameter W61TO61 = 0;
parameter W61TO62 = 0;
parameter W61TO63 = 0;
parameter W61TO64 = 0;
parameter W61TO65 = 0;
parameter W61TO66 = 0;
parameter W61TO67 = 0;
parameter W61TO68 = 0;
parameter W61TO69 = 0;
parameter W61TO70 = 0;
parameter W61TO71 = 0;
parameter W61TO72 = 0;
parameter W61TO73 = 0;
parameter W61TO74 = 0;
parameter W61TO75 = 0;
parameter W61TO76 = 0;
parameter W61TO77 = 0;
parameter W61TO78 = 0;
parameter W61TO79 = 0;
parameter W61TO80 = 0;
parameter W61TO81 = 0;
parameter W61TO82 = 0;
parameter W61TO83 = 0;
parameter W61TO84 = 0;
parameter W61TO85 = 0;
parameter W61TO86 = 0;
parameter W61TO87 = 0;
parameter W61TO88 = 0;
parameter W61TO89 = 0;
parameter W61TO90 = 0;
parameter W61TO91 = 0;
parameter W61TO92 = 0;
parameter W61TO93 = 0;
parameter W61TO94 = 0;
parameter W61TO95 = 0;
parameter W61TO96 = 0;
parameter W61TO97 = 0;
parameter W61TO98 = 0;
parameter W61TO99 = 0;
parameter W62TO0 = 0;
parameter W62TO1 = 0;
parameter W62TO2 = 0;
parameter W62TO3 = 0;
parameter W62TO4 = 0;
parameter W62TO5 = 0;
parameter W62TO6 = 0;
parameter W62TO7 = 0;
parameter W62TO8 = 0;
parameter W62TO9 = 0;
parameter W62TO10 = 0;
parameter W62TO11 = 0;
parameter W62TO12 = 0;
parameter W62TO13 = 0;
parameter W62TO14 = 0;
parameter W62TO15 = 0;
parameter W62TO16 = 0;
parameter W62TO17 = 0;
parameter W62TO18 = 0;
parameter W62TO19 = 0;
parameter W62TO20 = 0;
parameter W62TO21 = 0;
parameter W62TO22 = 0;
parameter W62TO23 = 0;
parameter W62TO24 = 0;
parameter W62TO25 = 0;
parameter W62TO26 = 0;
parameter W62TO27 = 0;
parameter W62TO28 = 0;
parameter W62TO29 = 0;
parameter W62TO30 = 0;
parameter W62TO31 = 0;
parameter W62TO32 = 0;
parameter W62TO33 = 0;
parameter W62TO34 = 0;
parameter W62TO35 = 0;
parameter W62TO36 = 0;
parameter W62TO37 = 0;
parameter W62TO38 = 0;
parameter W62TO39 = 0;
parameter W62TO40 = 0;
parameter W62TO41 = 0;
parameter W62TO42 = 0;
parameter W62TO43 = 0;
parameter W62TO44 = 0;
parameter W62TO45 = 0;
parameter W62TO46 = 0;
parameter W62TO47 = 0;
parameter W62TO48 = 0;
parameter W62TO49 = 0;
parameter W62TO50 = 0;
parameter W62TO51 = 0;
parameter W62TO52 = 0;
parameter W62TO53 = 0;
parameter W62TO54 = 0;
parameter W62TO55 = 0;
parameter W62TO56 = 0;
parameter W62TO57 = 0;
parameter W62TO58 = 0;
parameter W62TO59 = 0;
parameter W62TO60 = 0;
parameter W62TO61 = 0;
parameter W62TO62 = 0;
parameter W62TO63 = 0;
parameter W62TO64 = 0;
parameter W62TO65 = 0;
parameter W62TO66 = 0;
parameter W62TO67 = 0;
parameter W62TO68 = 0;
parameter W62TO69 = 0;
parameter W62TO70 = 0;
parameter W62TO71 = 0;
parameter W62TO72 = 0;
parameter W62TO73 = 0;
parameter W62TO74 = 0;
parameter W62TO75 = 0;
parameter W62TO76 = 0;
parameter W62TO77 = 0;
parameter W62TO78 = 0;
parameter W62TO79 = 0;
parameter W62TO80 = 0;
parameter W62TO81 = 0;
parameter W62TO82 = 0;
parameter W62TO83 = 0;
parameter W62TO84 = 0;
parameter W62TO85 = 0;
parameter W62TO86 = 0;
parameter W62TO87 = 0;
parameter W62TO88 = 0;
parameter W62TO89 = 0;
parameter W62TO90 = 0;
parameter W62TO91 = 0;
parameter W62TO92 = 0;
parameter W62TO93 = 0;
parameter W62TO94 = 0;
parameter W62TO95 = 0;
parameter W62TO96 = 0;
parameter W62TO97 = 0;
parameter W62TO98 = 0;
parameter W62TO99 = 0;
parameter W63TO0 = 0;
parameter W63TO1 = 0;
parameter W63TO2 = 0;
parameter W63TO3 = 0;
parameter W63TO4 = 0;
parameter W63TO5 = 0;
parameter W63TO6 = 0;
parameter W63TO7 = 0;
parameter W63TO8 = 0;
parameter W63TO9 = 0;
parameter W63TO10 = 0;
parameter W63TO11 = 0;
parameter W63TO12 = 0;
parameter W63TO13 = 0;
parameter W63TO14 = 0;
parameter W63TO15 = 0;
parameter W63TO16 = 0;
parameter W63TO17 = 0;
parameter W63TO18 = 0;
parameter W63TO19 = 0;
parameter W63TO20 = 0;
parameter W63TO21 = 0;
parameter W63TO22 = 0;
parameter W63TO23 = 0;
parameter W63TO24 = 0;
parameter W63TO25 = 0;
parameter W63TO26 = 0;
parameter W63TO27 = 0;
parameter W63TO28 = 0;
parameter W63TO29 = 0;
parameter W63TO30 = 0;
parameter W63TO31 = 0;
parameter W63TO32 = 0;
parameter W63TO33 = 0;
parameter W63TO34 = 0;
parameter W63TO35 = 0;
parameter W63TO36 = 0;
parameter W63TO37 = 0;
parameter W63TO38 = 0;
parameter W63TO39 = 0;
parameter W63TO40 = 0;
parameter W63TO41 = 0;
parameter W63TO42 = 0;
parameter W63TO43 = 0;
parameter W63TO44 = 0;
parameter W63TO45 = 0;
parameter W63TO46 = 0;
parameter W63TO47 = 0;
parameter W63TO48 = 0;
parameter W63TO49 = 0;
parameter W63TO50 = 0;
parameter W63TO51 = 0;
parameter W63TO52 = 0;
parameter W63TO53 = 0;
parameter W63TO54 = 0;
parameter W63TO55 = 0;
parameter W63TO56 = 0;
parameter W63TO57 = 0;
parameter W63TO58 = 0;
parameter W63TO59 = 0;
parameter W63TO60 = 0;
parameter W63TO61 = 0;
parameter W63TO62 = 0;
parameter W63TO63 = 0;
parameter W63TO64 = 0;
parameter W63TO65 = 0;
parameter W63TO66 = 0;
parameter W63TO67 = 0;
parameter W63TO68 = 0;
parameter W63TO69 = 0;
parameter W63TO70 = 0;
parameter W63TO71 = 0;
parameter W63TO72 = 0;
parameter W63TO73 = 0;
parameter W63TO74 = 0;
parameter W63TO75 = 0;
parameter W63TO76 = 0;
parameter W63TO77 = 0;
parameter W63TO78 = 0;
parameter W63TO79 = 0;
parameter W63TO80 = 0;
parameter W63TO81 = 0;
parameter W63TO82 = 0;
parameter W63TO83 = 0;
parameter W63TO84 = 0;
parameter W63TO85 = 0;
parameter W63TO86 = 0;
parameter W63TO87 = 0;
parameter W63TO88 = 0;
parameter W63TO89 = 0;
parameter W63TO90 = 0;
parameter W63TO91 = 0;
parameter W63TO92 = 0;
parameter W63TO93 = 0;
parameter W63TO94 = 0;
parameter W63TO95 = 0;
parameter W63TO96 = 0;
parameter W63TO97 = 0;
parameter W63TO98 = 0;
parameter W63TO99 = 0;

input wire clk;
input wire rst;

input signed [15:0] in0;
input signed [15:0] in1;
input signed [15:0] in2;
input signed [15:0] in3;
input signed [15:0] in4;
input signed [15:0] in5;
input signed [15:0] in6;
input signed [15:0] in7;
input signed [15:0] in8;
input signed [15:0] in9;
input signed [15:0] in10;
input signed [15:0] in11;
input signed [15:0] in12;
input signed [15:0] in13;
input signed [15:0] in14;
input signed [15:0] in15;
input signed [15:0] in16;
input signed [15:0] in17;
input signed [15:0] in18;
input signed [15:0] in19;
input signed [15:0] in20;
input signed [15:0] in21;
input signed [15:0] in22;
input signed [15:0] in23;
input signed [15:0] in24;
input signed [15:0] in25;
input signed [15:0] in26;
input signed [15:0] in27;
input signed [15:0] in28;
input signed [15:0] in29;
input signed [15:0] in30;
input signed [15:0] in31;
input signed [15:0] in32;
input signed [15:0] in33;
input signed [15:0] in34;
input signed [15:0] in35;
input signed [15:0] in36;
input signed [15:0] in37;
input signed [15:0] in38;
input signed [15:0] in39;
input signed [15:0] in40;
input signed [15:0] in41;
input signed [15:0] in42;
input signed [15:0] in43;
input signed [15:0] in44;
input signed [15:0] in45;
input signed [15:0] in46;
input signed [15:0] in47;
input signed [15:0] in48;
input signed [15:0] in49;
input signed [15:0] in50;
input signed [15:0] in51;
input signed [15:0] in52;
input signed [15:0] in53;
input signed [15:0] in54;
input signed [15:0] in55;
input signed [15:0] in56;
input signed [15:0] in57;
input signed [15:0] in58;
input signed [15:0] in59;
input signed [15:0] in60;
input signed [15:0] in61;
input signed [15:0] in62;
input signed [15:0] in63;

output signed [15:0] out0;
output signed [15:0] out1;
output signed [15:0] out2;
output signed [15:0] out3;
output signed [15:0] out4;
output signed [15:0] out5;
output signed [15:0] out6;
output signed [15:0] out7;
output signed [15:0] out8;
output signed [15:0] out9;
output signed [15:0] out10;
output signed [15:0] out11;
output signed [15:0] out12;
output signed [15:0] out13;
output signed [15:0] out14;
output signed [15:0] out15;
output signed [15:0] out16;
output signed [15:0] out17;
output signed [15:0] out18;
output signed [15:0] out19;
output signed [15:0] out20;
output signed [15:0] out21;
output signed [15:0] out22;
output signed [15:0] out23;
output signed [15:0] out24;
output signed [15:0] out25;
output signed [15:0] out26;
output signed [15:0] out27;
output signed [15:0] out28;
output signed [15:0] out29;
output signed [15:0] out30;
output signed [15:0] out31;
output signed [15:0] out32;
output signed [15:0] out33;
output signed [15:0] out34;
output signed [15:0] out35;
output signed [15:0] out36;
output signed [15:0] out37;
output signed [15:0] out38;
output signed [15:0] out39;
output signed [15:0] out40;
output signed [15:0] out41;
output signed [15:0] out42;
output signed [15:0] out43;
output signed [15:0] out44;
output signed [15:0] out45;
output signed [15:0] out46;
output signed [15:0] out47;
output signed [15:0] out48;
output signed [15:0] out49;
output signed [15:0] out50;
output signed [15:0] out51;
output signed [15:0] out52;
output signed [15:0] out53;
output signed [15:0] out54;
output signed [15:0] out55;
output signed [15:0] out56;
output signed [15:0] out57;
output signed [15:0] out58;
output signed [15:0] out59;
output signed [15:0] out60;
output signed [15:0] out61;
output signed [15:0] out62;
output signed [15:0] out63;
output signed [15:0] out64;
output signed [15:0] out65;
output signed [15:0] out66;
output signed [15:0] out67;
output signed [15:0] out68;
output signed [15:0] out69;
output signed [15:0] out70;
output signed [15:0] out71;
output signed [15:0] out72;
output signed [15:0] out73;
output signed [15:0] out74;
output signed [15:0] out75;
output signed [15:0] out76;
output signed [15:0] out77;
output signed [15:0] out78;
output signed [15:0] out79;
output signed [15:0] out80;
output signed [15:0] out81;
output signed [15:0] out82;
output signed [15:0] out83;
output signed [15:0] out84;
output signed [15:0] out85;
output signed [15:0] out86;
output signed [15:0] out87;
output signed [15:0] out88;
output signed [15:0] out89;
output signed [15:0] out90;
output signed [15:0] out91;
output signed [15:0] out92;
output signed [15:0] out93;
output signed [15:0] out94;
output signed [15:0] out95;
output signed [15:0] out96;
output signed [15:0] out97;
output signed [15:0] out98;
output signed [15:0] out99;

neuron64in #(.W0(W0TO0), .W1(W1TO0), .W2(W2TO0), .W3(W3TO0), .W4(W4TO0), .W5(W5TO0), .W6(W6TO0), .W7(W7TO0), .W8(W8TO0), .W9(W9TO0), .W10(W10TO0), .W11(W11TO0), .W12(W12TO0), .W13(W13TO0), .W14(W14TO0), .W15(W15TO0), .W16(W16TO0), .W17(W17TO0), .W18(W18TO0), .W19(W19TO0), .W20(W20TO0), .W21(W21TO0), .W22(W22TO0), .W23(W23TO0), .W24(W24TO0), .W25(W25TO0), .W26(W26TO0), .W27(W27TO0), .W28(W28TO0), .W29(W29TO0), .W30(W30TO0), .W31(W31TO0), .W32(W32TO0), .W33(W33TO0), .W34(W34TO0), .W35(W35TO0), .W36(W36TO0), .W37(W37TO0), .W38(W38TO0), .W39(W39TO0), .W40(W40TO0), .W41(W41TO0), .W42(W42TO0), .W43(W43TO0), .W44(W44TO0), .W45(W45TO0), .W46(W46TO0), .W47(W47TO0), .W48(W48TO0), .W49(W49TO0), .W50(W50TO0), .W51(W51TO0), .W52(W52TO0), .W53(W53TO0), .W54(W54TO0), .W55(W55TO0), .W56(W56TO0), .W57(W57TO0), .W58(W58TO0), .W59(W59TO0), .W60(W60TO0), .W61(W61TO0), .W62(W62TO0), .W63(W63TO0)) neuron0(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out0));
neuron64in #(.W0(W0TO1), .W1(W1TO1), .W2(W2TO1), .W3(W3TO1), .W4(W4TO1), .W5(W5TO1), .W6(W6TO1), .W7(W7TO1), .W8(W8TO1), .W9(W9TO1), .W10(W10TO1), .W11(W11TO1), .W12(W12TO1), .W13(W13TO1), .W14(W14TO1), .W15(W15TO1), .W16(W16TO1), .W17(W17TO1), .W18(W18TO1), .W19(W19TO1), .W20(W20TO1), .W21(W21TO1), .W22(W22TO1), .W23(W23TO1), .W24(W24TO1), .W25(W25TO1), .W26(W26TO1), .W27(W27TO1), .W28(W28TO1), .W29(W29TO1), .W30(W30TO1), .W31(W31TO1), .W32(W32TO1), .W33(W33TO1), .W34(W34TO1), .W35(W35TO1), .W36(W36TO1), .W37(W37TO1), .W38(W38TO1), .W39(W39TO1), .W40(W40TO1), .W41(W41TO1), .W42(W42TO1), .W43(W43TO1), .W44(W44TO1), .W45(W45TO1), .W46(W46TO1), .W47(W47TO1), .W48(W48TO1), .W49(W49TO1), .W50(W50TO1), .W51(W51TO1), .W52(W52TO1), .W53(W53TO1), .W54(W54TO1), .W55(W55TO1), .W56(W56TO1), .W57(W57TO1), .W58(W58TO1), .W59(W59TO1), .W60(W60TO1), .W61(W61TO1), .W62(W62TO1), .W63(W63TO1)) neuron1(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out1));
neuron64in #(.W0(W0TO2), .W1(W1TO2), .W2(W2TO2), .W3(W3TO2), .W4(W4TO2), .W5(W5TO2), .W6(W6TO2), .W7(W7TO2), .W8(W8TO2), .W9(W9TO2), .W10(W10TO2), .W11(W11TO2), .W12(W12TO2), .W13(W13TO2), .W14(W14TO2), .W15(W15TO2), .W16(W16TO2), .W17(W17TO2), .W18(W18TO2), .W19(W19TO2), .W20(W20TO2), .W21(W21TO2), .W22(W22TO2), .W23(W23TO2), .W24(W24TO2), .W25(W25TO2), .W26(W26TO2), .W27(W27TO2), .W28(W28TO2), .W29(W29TO2), .W30(W30TO2), .W31(W31TO2), .W32(W32TO2), .W33(W33TO2), .W34(W34TO2), .W35(W35TO2), .W36(W36TO2), .W37(W37TO2), .W38(W38TO2), .W39(W39TO2), .W40(W40TO2), .W41(W41TO2), .W42(W42TO2), .W43(W43TO2), .W44(W44TO2), .W45(W45TO2), .W46(W46TO2), .W47(W47TO2), .W48(W48TO2), .W49(W49TO2), .W50(W50TO2), .W51(W51TO2), .W52(W52TO2), .W53(W53TO2), .W54(W54TO2), .W55(W55TO2), .W56(W56TO2), .W57(W57TO2), .W58(W58TO2), .W59(W59TO2), .W60(W60TO2), .W61(W61TO2), .W62(W62TO2), .W63(W63TO2)) neuron2(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out2));
neuron64in #(.W0(W0TO3), .W1(W1TO3), .W2(W2TO3), .W3(W3TO3), .W4(W4TO3), .W5(W5TO3), .W6(W6TO3), .W7(W7TO3), .W8(W8TO3), .W9(W9TO3), .W10(W10TO3), .W11(W11TO3), .W12(W12TO3), .W13(W13TO3), .W14(W14TO3), .W15(W15TO3), .W16(W16TO3), .W17(W17TO3), .W18(W18TO3), .W19(W19TO3), .W20(W20TO3), .W21(W21TO3), .W22(W22TO3), .W23(W23TO3), .W24(W24TO3), .W25(W25TO3), .W26(W26TO3), .W27(W27TO3), .W28(W28TO3), .W29(W29TO3), .W30(W30TO3), .W31(W31TO3), .W32(W32TO3), .W33(W33TO3), .W34(W34TO3), .W35(W35TO3), .W36(W36TO3), .W37(W37TO3), .W38(W38TO3), .W39(W39TO3), .W40(W40TO3), .W41(W41TO3), .W42(W42TO3), .W43(W43TO3), .W44(W44TO3), .W45(W45TO3), .W46(W46TO3), .W47(W47TO3), .W48(W48TO3), .W49(W49TO3), .W50(W50TO3), .W51(W51TO3), .W52(W52TO3), .W53(W53TO3), .W54(W54TO3), .W55(W55TO3), .W56(W56TO3), .W57(W57TO3), .W58(W58TO3), .W59(W59TO3), .W60(W60TO3), .W61(W61TO3), .W62(W62TO3), .W63(W63TO3)) neuron3(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out3));
neuron64in #(.W0(W0TO4), .W1(W1TO4), .W2(W2TO4), .W3(W3TO4), .W4(W4TO4), .W5(W5TO4), .W6(W6TO4), .W7(W7TO4), .W8(W8TO4), .W9(W9TO4), .W10(W10TO4), .W11(W11TO4), .W12(W12TO4), .W13(W13TO4), .W14(W14TO4), .W15(W15TO4), .W16(W16TO4), .W17(W17TO4), .W18(W18TO4), .W19(W19TO4), .W20(W20TO4), .W21(W21TO4), .W22(W22TO4), .W23(W23TO4), .W24(W24TO4), .W25(W25TO4), .W26(W26TO4), .W27(W27TO4), .W28(W28TO4), .W29(W29TO4), .W30(W30TO4), .W31(W31TO4), .W32(W32TO4), .W33(W33TO4), .W34(W34TO4), .W35(W35TO4), .W36(W36TO4), .W37(W37TO4), .W38(W38TO4), .W39(W39TO4), .W40(W40TO4), .W41(W41TO4), .W42(W42TO4), .W43(W43TO4), .W44(W44TO4), .W45(W45TO4), .W46(W46TO4), .W47(W47TO4), .W48(W48TO4), .W49(W49TO4), .W50(W50TO4), .W51(W51TO4), .W52(W52TO4), .W53(W53TO4), .W54(W54TO4), .W55(W55TO4), .W56(W56TO4), .W57(W57TO4), .W58(W58TO4), .W59(W59TO4), .W60(W60TO4), .W61(W61TO4), .W62(W62TO4), .W63(W63TO4)) neuron4(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out4));
neuron64in #(.W0(W0TO5), .W1(W1TO5), .W2(W2TO5), .W3(W3TO5), .W4(W4TO5), .W5(W5TO5), .W6(W6TO5), .W7(W7TO5), .W8(W8TO5), .W9(W9TO5), .W10(W10TO5), .W11(W11TO5), .W12(W12TO5), .W13(W13TO5), .W14(W14TO5), .W15(W15TO5), .W16(W16TO5), .W17(W17TO5), .W18(W18TO5), .W19(W19TO5), .W20(W20TO5), .W21(W21TO5), .W22(W22TO5), .W23(W23TO5), .W24(W24TO5), .W25(W25TO5), .W26(W26TO5), .W27(W27TO5), .W28(W28TO5), .W29(W29TO5), .W30(W30TO5), .W31(W31TO5), .W32(W32TO5), .W33(W33TO5), .W34(W34TO5), .W35(W35TO5), .W36(W36TO5), .W37(W37TO5), .W38(W38TO5), .W39(W39TO5), .W40(W40TO5), .W41(W41TO5), .W42(W42TO5), .W43(W43TO5), .W44(W44TO5), .W45(W45TO5), .W46(W46TO5), .W47(W47TO5), .W48(W48TO5), .W49(W49TO5), .W50(W50TO5), .W51(W51TO5), .W52(W52TO5), .W53(W53TO5), .W54(W54TO5), .W55(W55TO5), .W56(W56TO5), .W57(W57TO5), .W58(W58TO5), .W59(W59TO5), .W60(W60TO5), .W61(W61TO5), .W62(W62TO5), .W63(W63TO5)) neuron5(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out5));
neuron64in #(.W0(W0TO6), .W1(W1TO6), .W2(W2TO6), .W3(W3TO6), .W4(W4TO6), .W5(W5TO6), .W6(W6TO6), .W7(W7TO6), .W8(W8TO6), .W9(W9TO6), .W10(W10TO6), .W11(W11TO6), .W12(W12TO6), .W13(W13TO6), .W14(W14TO6), .W15(W15TO6), .W16(W16TO6), .W17(W17TO6), .W18(W18TO6), .W19(W19TO6), .W20(W20TO6), .W21(W21TO6), .W22(W22TO6), .W23(W23TO6), .W24(W24TO6), .W25(W25TO6), .W26(W26TO6), .W27(W27TO6), .W28(W28TO6), .W29(W29TO6), .W30(W30TO6), .W31(W31TO6), .W32(W32TO6), .W33(W33TO6), .W34(W34TO6), .W35(W35TO6), .W36(W36TO6), .W37(W37TO6), .W38(W38TO6), .W39(W39TO6), .W40(W40TO6), .W41(W41TO6), .W42(W42TO6), .W43(W43TO6), .W44(W44TO6), .W45(W45TO6), .W46(W46TO6), .W47(W47TO6), .W48(W48TO6), .W49(W49TO6), .W50(W50TO6), .W51(W51TO6), .W52(W52TO6), .W53(W53TO6), .W54(W54TO6), .W55(W55TO6), .W56(W56TO6), .W57(W57TO6), .W58(W58TO6), .W59(W59TO6), .W60(W60TO6), .W61(W61TO6), .W62(W62TO6), .W63(W63TO6)) neuron6(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out6));
neuron64in #(.W0(W0TO7), .W1(W1TO7), .W2(W2TO7), .W3(W3TO7), .W4(W4TO7), .W5(W5TO7), .W6(W6TO7), .W7(W7TO7), .W8(W8TO7), .W9(W9TO7), .W10(W10TO7), .W11(W11TO7), .W12(W12TO7), .W13(W13TO7), .W14(W14TO7), .W15(W15TO7), .W16(W16TO7), .W17(W17TO7), .W18(W18TO7), .W19(W19TO7), .W20(W20TO7), .W21(W21TO7), .W22(W22TO7), .W23(W23TO7), .W24(W24TO7), .W25(W25TO7), .W26(W26TO7), .W27(W27TO7), .W28(W28TO7), .W29(W29TO7), .W30(W30TO7), .W31(W31TO7), .W32(W32TO7), .W33(W33TO7), .W34(W34TO7), .W35(W35TO7), .W36(W36TO7), .W37(W37TO7), .W38(W38TO7), .W39(W39TO7), .W40(W40TO7), .W41(W41TO7), .W42(W42TO7), .W43(W43TO7), .W44(W44TO7), .W45(W45TO7), .W46(W46TO7), .W47(W47TO7), .W48(W48TO7), .W49(W49TO7), .W50(W50TO7), .W51(W51TO7), .W52(W52TO7), .W53(W53TO7), .W54(W54TO7), .W55(W55TO7), .W56(W56TO7), .W57(W57TO7), .W58(W58TO7), .W59(W59TO7), .W60(W60TO7), .W61(W61TO7), .W62(W62TO7), .W63(W63TO7)) neuron7(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out7));
neuron64in #(.W0(W0TO8), .W1(W1TO8), .W2(W2TO8), .W3(W3TO8), .W4(W4TO8), .W5(W5TO8), .W6(W6TO8), .W7(W7TO8), .W8(W8TO8), .W9(W9TO8), .W10(W10TO8), .W11(W11TO8), .W12(W12TO8), .W13(W13TO8), .W14(W14TO8), .W15(W15TO8), .W16(W16TO8), .W17(W17TO8), .W18(W18TO8), .W19(W19TO8), .W20(W20TO8), .W21(W21TO8), .W22(W22TO8), .W23(W23TO8), .W24(W24TO8), .W25(W25TO8), .W26(W26TO8), .W27(W27TO8), .W28(W28TO8), .W29(W29TO8), .W30(W30TO8), .W31(W31TO8), .W32(W32TO8), .W33(W33TO8), .W34(W34TO8), .W35(W35TO8), .W36(W36TO8), .W37(W37TO8), .W38(W38TO8), .W39(W39TO8), .W40(W40TO8), .W41(W41TO8), .W42(W42TO8), .W43(W43TO8), .W44(W44TO8), .W45(W45TO8), .W46(W46TO8), .W47(W47TO8), .W48(W48TO8), .W49(W49TO8), .W50(W50TO8), .W51(W51TO8), .W52(W52TO8), .W53(W53TO8), .W54(W54TO8), .W55(W55TO8), .W56(W56TO8), .W57(W57TO8), .W58(W58TO8), .W59(W59TO8), .W60(W60TO8), .W61(W61TO8), .W62(W62TO8), .W63(W63TO8)) neuron8(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out8));
neuron64in #(.W0(W0TO9), .W1(W1TO9), .W2(W2TO9), .W3(W3TO9), .W4(W4TO9), .W5(W5TO9), .W6(W6TO9), .W7(W7TO9), .W8(W8TO9), .W9(W9TO9), .W10(W10TO9), .W11(W11TO9), .W12(W12TO9), .W13(W13TO9), .W14(W14TO9), .W15(W15TO9), .W16(W16TO9), .W17(W17TO9), .W18(W18TO9), .W19(W19TO9), .W20(W20TO9), .W21(W21TO9), .W22(W22TO9), .W23(W23TO9), .W24(W24TO9), .W25(W25TO9), .W26(W26TO9), .W27(W27TO9), .W28(W28TO9), .W29(W29TO9), .W30(W30TO9), .W31(W31TO9), .W32(W32TO9), .W33(W33TO9), .W34(W34TO9), .W35(W35TO9), .W36(W36TO9), .W37(W37TO9), .W38(W38TO9), .W39(W39TO9), .W40(W40TO9), .W41(W41TO9), .W42(W42TO9), .W43(W43TO9), .W44(W44TO9), .W45(W45TO9), .W46(W46TO9), .W47(W47TO9), .W48(W48TO9), .W49(W49TO9), .W50(W50TO9), .W51(W51TO9), .W52(W52TO9), .W53(W53TO9), .W54(W54TO9), .W55(W55TO9), .W56(W56TO9), .W57(W57TO9), .W58(W58TO9), .W59(W59TO9), .W60(W60TO9), .W61(W61TO9), .W62(W62TO9), .W63(W63TO9)) neuron9(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out9));
neuron64in #(.W0(W0TO10), .W1(W1TO10), .W2(W2TO10), .W3(W3TO10), .W4(W4TO10), .W5(W5TO10), .W6(W6TO10), .W7(W7TO10), .W8(W8TO10), .W9(W9TO10), .W10(W10TO10), .W11(W11TO10), .W12(W12TO10), .W13(W13TO10), .W14(W14TO10), .W15(W15TO10), .W16(W16TO10), .W17(W17TO10), .W18(W18TO10), .W19(W19TO10), .W20(W20TO10), .W21(W21TO10), .W22(W22TO10), .W23(W23TO10), .W24(W24TO10), .W25(W25TO10), .W26(W26TO10), .W27(W27TO10), .W28(W28TO10), .W29(W29TO10), .W30(W30TO10), .W31(W31TO10), .W32(W32TO10), .W33(W33TO10), .W34(W34TO10), .W35(W35TO10), .W36(W36TO10), .W37(W37TO10), .W38(W38TO10), .W39(W39TO10), .W40(W40TO10), .W41(W41TO10), .W42(W42TO10), .W43(W43TO10), .W44(W44TO10), .W45(W45TO10), .W46(W46TO10), .W47(W47TO10), .W48(W48TO10), .W49(W49TO10), .W50(W50TO10), .W51(W51TO10), .W52(W52TO10), .W53(W53TO10), .W54(W54TO10), .W55(W55TO10), .W56(W56TO10), .W57(W57TO10), .W58(W58TO10), .W59(W59TO10), .W60(W60TO10), .W61(W61TO10), .W62(W62TO10), .W63(W63TO10)) neuron10(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out10));
neuron64in #(.W0(W0TO11), .W1(W1TO11), .W2(W2TO11), .W3(W3TO11), .W4(W4TO11), .W5(W5TO11), .W6(W6TO11), .W7(W7TO11), .W8(W8TO11), .W9(W9TO11), .W10(W10TO11), .W11(W11TO11), .W12(W12TO11), .W13(W13TO11), .W14(W14TO11), .W15(W15TO11), .W16(W16TO11), .W17(W17TO11), .W18(W18TO11), .W19(W19TO11), .W20(W20TO11), .W21(W21TO11), .W22(W22TO11), .W23(W23TO11), .W24(W24TO11), .W25(W25TO11), .W26(W26TO11), .W27(W27TO11), .W28(W28TO11), .W29(W29TO11), .W30(W30TO11), .W31(W31TO11), .W32(W32TO11), .W33(W33TO11), .W34(W34TO11), .W35(W35TO11), .W36(W36TO11), .W37(W37TO11), .W38(W38TO11), .W39(W39TO11), .W40(W40TO11), .W41(W41TO11), .W42(W42TO11), .W43(W43TO11), .W44(W44TO11), .W45(W45TO11), .W46(W46TO11), .W47(W47TO11), .W48(W48TO11), .W49(W49TO11), .W50(W50TO11), .W51(W51TO11), .W52(W52TO11), .W53(W53TO11), .W54(W54TO11), .W55(W55TO11), .W56(W56TO11), .W57(W57TO11), .W58(W58TO11), .W59(W59TO11), .W60(W60TO11), .W61(W61TO11), .W62(W62TO11), .W63(W63TO11)) neuron11(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out11));
neuron64in #(.W0(W0TO12), .W1(W1TO12), .W2(W2TO12), .W3(W3TO12), .W4(W4TO12), .W5(W5TO12), .W6(W6TO12), .W7(W7TO12), .W8(W8TO12), .W9(W9TO12), .W10(W10TO12), .W11(W11TO12), .W12(W12TO12), .W13(W13TO12), .W14(W14TO12), .W15(W15TO12), .W16(W16TO12), .W17(W17TO12), .W18(W18TO12), .W19(W19TO12), .W20(W20TO12), .W21(W21TO12), .W22(W22TO12), .W23(W23TO12), .W24(W24TO12), .W25(W25TO12), .W26(W26TO12), .W27(W27TO12), .W28(W28TO12), .W29(W29TO12), .W30(W30TO12), .W31(W31TO12), .W32(W32TO12), .W33(W33TO12), .W34(W34TO12), .W35(W35TO12), .W36(W36TO12), .W37(W37TO12), .W38(W38TO12), .W39(W39TO12), .W40(W40TO12), .W41(W41TO12), .W42(W42TO12), .W43(W43TO12), .W44(W44TO12), .W45(W45TO12), .W46(W46TO12), .W47(W47TO12), .W48(W48TO12), .W49(W49TO12), .W50(W50TO12), .W51(W51TO12), .W52(W52TO12), .W53(W53TO12), .W54(W54TO12), .W55(W55TO12), .W56(W56TO12), .W57(W57TO12), .W58(W58TO12), .W59(W59TO12), .W60(W60TO12), .W61(W61TO12), .W62(W62TO12), .W63(W63TO12)) neuron12(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out12));
neuron64in #(.W0(W0TO13), .W1(W1TO13), .W2(W2TO13), .W3(W3TO13), .W4(W4TO13), .W5(W5TO13), .W6(W6TO13), .W7(W7TO13), .W8(W8TO13), .W9(W9TO13), .W10(W10TO13), .W11(W11TO13), .W12(W12TO13), .W13(W13TO13), .W14(W14TO13), .W15(W15TO13), .W16(W16TO13), .W17(W17TO13), .W18(W18TO13), .W19(W19TO13), .W20(W20TO13), .W21(W21TO13), .W22(W22TO13), .W23(W23TO13), .W24(W24TO13), .W25(W25TO13), .W26(W26TO13), .W27(W27TO13), .W28(W28TO13), .W29(W29TO13), .W30(W30TO13), .W31(W31TO13), .W32(W32TO13), .W33(W33TO13), .W34(W34TO13), .W35(W35TO13), .W36(W36TO13), .W37(W37TO13), .W38(W38TO13), .W39(W39TO13), .W40(W40TO13), .W41(W41TO13), .W42(W42TO13), .W43(W43TO13), .W44(W44TO13), .W45(W45TO13), .W46(W46TO13), .W47(W47TO13), .W48(W48TO13), .W49(W49TO13), .W50(W50TO13), .W51(W51TO13), .W52(W52TO13), .W53(W53TO13), .W54(W54TO13), .W55(W55TO13), .W56(W56TO13), .W57(W57TO13), .W58(W58TO13), .W59(W59TO13), .W60(W60TO13), .W61(W61TO13), .W62(W62TO13), .W63(W63TO13)) neuron13(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out13));
neuron64in #(.W0(W0TO14), .W1(W1TO14), .W2(W2TO14), .W3(W3TO14), .W4(W4TO14), .W5(W5TO14), .W6(W6TO14), .W7(W7TO14), .W8(W8TO14), .W9(W9TO14), .W10(W10TO14), .W11(W11TO14), .W12(W12TO14), .W13(W13TO14), .W14(W14TO14), .W15(W15TO14), .W16(W16TO14), .W17(W17TO14), .W18(W18TO14), .W19(W19TO14), .W20(W20TO14), .W21(W21TO14), .W22(W22TO14), .W23(W23TO14), .W24(W24TO14), .W25(W25TO14), .W26(W26TO14), .W27(W27TO14), .W28(W28TO14), .W29(W29TO14), .W30(W30TO14), .W31(W31TO14), .W32(W32TO14), .W33(W33TO14), .W34(W34TO14), .W35(W35TO14), .W36(W36TO14), .W37(W37TO14), .W38(W38TO14), .W39(W39TO14), .W40(W40TO14), .W41(W41TO14), .W42(W42TO14), .W43(W43TO14), .W44(W44TO14), .W45(W45TO14), .W46(W46TO14), .W47(W47TO14), .W48(W48TO14), .W49(W49TO14), .W50(W50TO14), .W51(W51TO14), .W52(W52TO14), .W53(W53TO14), .W54(W54TO14), .W55(W55TO14), .W56(W56TO14), .W57(W57TO14), .W58(W58TO14), .W59(W59TO14), .W60(W60TO14), .W61(W61TO14), .W62(W62TO14), .W63(W63TO14)) neuron14(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out14));
neuron64in #(.W0(W0TO15), .W1(W1TO15), .W2(W2TO15), .W3(W3TO15), .W4(W4TO15), .W5(W5TO15), .W6(W6TO15), .W7(W7TO15), .W8(W8TO15), .W9(W9TO15), .W10(W10TO15), .W11(W11TO15), .W12(W12TO15), .W13(W13TO15), .W14(W14TO15), .W15(W15TO15), .W16(W16TO15), .W17(W17TO15), .W18(W18TO15), .W19(W19TO15), .W20(W20TO15), .W21(W21TO15), .W22(W22TO15), .W23(W23TO15), .W24(W24TO15), .W25(W25TO15), .W26(W26TO15), .W27(W27TO15), .W28(W28TO15), .W29(W29TO15), .W30(W30TO15), .W31(W31TO15), .W32(W32TO15), .W33(W33TO15), .W34(W34TO15), .W35(W35TO15), .W36(W36TO15), .W37(W37TO15), .W38(W38TO15), .W39(W39TO15), .W40(W40TO15), .W41(W41TO15), .W42(W42TO15), .W43(W43TO15), .W44(W44TO15), .W45(W45TO15), .W46(W46TO15), .W47(W47TO15), .W48(W48TO15), .W49(W49TO15), .W50(W50TO15), .W51(W51TO15), .W52(W52TO15), .W53(W53TO15), .W54(W54TO15), .W55(W55TO15), .W56(W56TO15), .W57(W57TO15), .W58(W58TO15), .W59(W59TO15), .W60(W60TO15), .W61(W61TO15), .W62(W62TO15), .W63(W63TO15)) neuron15(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out15));
neuron64in #(.W0(W0TO16), .W1(W1TO16), .W2(W2TO16), .W3(W3TO16), .W4(W4TO16), .W5(W5TO16), .W6(W6TO16), .W7(W7TO16), .W8(W8TO16), .W9(W9TO16), .W10(W10TO16), .W11(W11TO16), .W12(W12TO16), .W13(W13TO16), .W14(W14TO16), .W15(W15TO16), .W16(W16TO16), .W17(W17TO16), .W18(W18TO16), .W19(W19TO16), .W20(W20TO16), .W21(W21TO16), .W22(W22TO16), .W23(W23TO16), .W24(W24TO16), .W25(W25TO16), .W26(W26TO16), .W27(W27TO16), .W28(W28TO16), .W29(W29TO16), .W30(W30TO16), .W31(W31TO16), .W32(W32TO16), .W33(W33TO16), .W34(W34TO16), .W35(W35TO16), .W36(W36TO16), .W37(W37TO16), .W38(W38TO16), .W39(W39TO16), .W40(W40TO16), .W41(W41TO16), .W42(W42TO16), .W43(W43TO16), .W44(W44TO16), .W45(W45TO16), .W46(W46TO16), .W47(W47TO16), .W48(W48TO16), .W49(W49TO16), .W50(W50TO16), .W51(W51TO16), .W52(W52TO16), .W53(W53TO16), .W54(W54TO16), .W55(W55TO16), .W56(W56TO16), .W57(W57TO16), .W58(W58TO16), .W59(W59TO16), .W60(W60TO16), .W61(W61TO16), .W62(W62TO16), .W63(W63TO16)) neuron16(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out16));
neuron64in #(.W0(W0TO17), .W1(W1TO17), .W2(W2TO17), .W3(W3TO17), .W4(W4TO17), .W5(W5TO17), .W6(W6TO17), .W7(W7TO17), .W8(W8TO17), .W9(W9TO17), .W10(W10TO17), .W11(W11TO17), .W12(W12TO17), .W13(W13TO17), .W14(W14TO17), .W15(W15TO17), .W16(W16TO17), .W17(W17TO17), .W18(W18TO17), .W19(W19TO17), .W20(W20TO17), .W21(W21TO17), .W22(W22TO17), .W23(W23TO17), .W24(W24TO17), .W25(W25TO17), .W26(W26TO17), .W27(W27TO17), .W28(W28TO17), .W29(W29TO17), .W30(W30TO17), .W31(W31TO17), .W32(W32TO17), .W33(W33TO17), .W34(W34TO17), .W35(W35TO17), .W36(W36TO17), .W37(W37TO17), .W38(W38TO17), .W39(W39TO17), .W40(W40TO17), .W41(W41TO17), .W42(W42TO17), .W43(W43TO17), .W44(W44TO17), .W45(W45TO17), .W46(W46TO17), .W47(W47TO17), .W48(W48TO17), .W49(W49TO17), .W50(W50TO17), .W51(W51TO17), .W52(W52TO17), .W53(W53TO17), .W54(W54TO17), .W55(W55TO17), .W56(W56TO17), .W57(W57TO17), .W58(W58TO17), .W59(W59TO17), .W60(W60TO17), .W61(W61TO17), .W62(W62TO17), .W63(W63TO17)) neuron17(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out17));
neuron64in #(.W0(W0TO18), .W1(W1TO18), .W2(W2TO18), .W3(W3TO18), .W4(W4TO18), .W5(W5TO18), .W6(W6TO18), .W7(W7TO18), .W8(W8TO18), .W9(W9TO18), .W10(W10TO18), .W11(W11TO18), .W12(W12TO18), .W13(W13TO18), .W14(W14TO18), .W15(W15TO18), .W16(W16TO18), .W17(W17TO18), .W18(W18TO18), .W19(W19TO18), .W20(W20TO18), .W21(W21TO18), .W22(W22TO18), .W23(W23TO18), .W24(W24TO18), .W25(W25TO18), .W26(W26TO18), .W27(W27TO18), .W28(W28TO18), .W29(W29TO18), .W30(W30TO18), .W31(W31TO18), .W32(W32TO18), .W33(W33TO18), .W34(W34TO18), .W35(W35TO18), .W36(W36TO18), .W37(W37TO18), .W38(W38TO18), .W39(W39TO18), .W40(W40TO18), .W41(W41TO18), .W42(W42TO18), .W43(W43TO18), .W44(W44TO18), .W45(W45TO18), .W46(W46TO18), .W47(W47TO18), .W48(W48TO18), .W49(W49TO18), .W50(W50TO18), .W51(W51TO18), .W52(W52TO18), .W53(W53TO18), .W54(W54TO18), .W55(W55TO18), .W56(W56TO18), .W57(W57TO18), .W58(W58TO18), .W59(W59TO18), .W60(W60TO18), .W61(W61TO18), .W62(W62TO18), .W63(W63TO18)) neuron18(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out18));
neuron64in #(.W0(W0TO19), .W1(W1TO19), .W2(W2TO19), .W3(W3TO19), .W4(W4TO19), .W5(W5TO19), .W6(W6TO19), .W7(W7TO19), .W8(W8TO19), .W9(W9TO19), .W10(W10TO19), .W11(W11TO19), .W12(W12TO19), .W13(W13TO19), .W14(W14TO19), .W15(W15TO19), .W16(W16TO19), .W17(W17TO19), .W18(W18TO19), .W19(W19TO19), .W20(W20TO19), .W21(W21TO19), .W22(W22TO19), .W23(W23TO19), .W24(W24TO19), .W25(W25TO19), .W26(W26TO19), .W27(W27TO19), .W28(W28TO19), .W29(W29TO19), .W30(W30TO19), .W31(W31TO19), .W32(W32TO19), .W33(W33TO19), .W34(W34TO19), .W35(W35TO19), .W36(W36TO19), .W37(W37TO19), .W38(W38TO19), .W39(W39TO19), .W40(W40TO19), .W41(W41TO19), .W42(W42TO19), .W43(W43TO19), .W44(W44TO19), .W45(W45TO19), .W46(W46TO19), .W47(W47TO19), .W48(W48TO19), .W49(W49TO19), .W50(W50TO19), .W51(W51TO19), .W52(W52TO19), .W53(W53TO19), .W54(W54TO19), .W55(W55TO19), .W56(W56TO19), .W57(W57TO19), .W58(W58TO19), .W59(W59TO19), .W60(W60TO19), .W61(W61TO19), .W62(W62TO19), .W63(W63TO19)) neuron19(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out19));
neuron64in #(.W0(W0TO20), .W1(W1TO20), .W2(W2TO20), .W3(W3TO20), .W4(W4TO20), .W5(W5TO20), .W6(W6TO20), .W7(W7TO20), .W8(W8TO20), .W9(W9TO20), .W10(W10TO20), .W11(W11TO20), .W12(W12TO20), .W13(W13TO20), .W14(W14TO20), .W15(W15TO20), .W16(W16TO20), .W17(W17TO20), .W18(W18TO20), .W19(W19TO20), .W20(W20TO20), .W21(W21TO20), .W22(W22TO20), .W23(W23TO20), .W24(W24TO20), .W25(W25TO20), .W26(W26TO20), .W27(W27TO20), .W28(W28TO20), .W29(W29TO20), .W30(W30TO20), .W31(W31TO20), .W32(W32TO20), .W33(W33TO20), .W34(W34TO20), .W35(W35TO20), .W36(W36TO20), .W37(W37TO20), .W38(W38TO20), .W39(W39TO20), .W40(W40TO20), .W41(W41TO20), .W42(W42TO20), .W43(W43TO20), .W44(W44TO20), .W45(W45TO20), .W46(W46TO20), .W47(W47TO20), .W48(W48TO20), .W49(W49TO20), .W50(W50TO20), .W51(W51TO20), .W52(W52TO20), .W53(W53TO20), .W54(W54TO20), .W55(W55TO20), .W56(W56TO20), .W57(W57TO20), .W58(W58TO20), .W59(W59TO20), .W60(W60TO20), .W61(W61TO20), .W62(W62TO20), .W63(W63TO20)) neuron20(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out20));
neuron64in #(.W0(W0TO21), .W1(W1TO21), .W2(W2TO21), .W3(W3TO21), .W4(W4TO21), .W5(W5TO21), .W6(W6TO21), .W7(W7TO21), .W8(W8TO21), .W9(W9TO21), .W10(W10TO21), .W11(W11TO21), .W12(W12TO21), .W13(W13TO21), .W14(W14TO21), .W15(W15TO21), .W16(W16TO21), .W17(W17TO21), .W18(W18TO21), .W19(W19TO21), .W20(W20TO21), .W21(W21TO21), .W22(W22TO21), .W23(W23TO21), .W24(W24TO21), .W25(W25TO21), .W26(W26TO21), .W27(W27TO21), .W28(W28TO21), .W29(W29TO21), .W30(W30TO21), .W31(W31TO21), .W32(W32TO21), .W33(W33TO21), .W34(W34TO21), .W35(W35TO21), .W36(W36TO21), .W37(W37TO21), .W38(W38TO21), .W39(W39TO21), .W40(W40TO21), .W41(W41TO21), .W42(W42TO21), .W43(W43TO21), .W44(W44TO21), .W45(W45TO21), .W46(W46TO21), .W47(W47TO21), .W48(W48TO21), .W49(W49TO21), .W50(W50TO21), .W51(W51TO21), .W52(W52TO21), .W53(W53TO21), .W54(W54TO21), .W55(W55TO21), .W56(W56TO21), .W57(W57TO21), .W58(W58TO21), .W59(W59TO21), .W60(W60TO21), .W61(W61TO21), .W62(W62TO21), .W63(W63TO21)) neuron21(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out21));
neuron64in #(.W0(W0TO22), .W1(W1TO22), .W2(W2TO22), .W3(W3TO22), .W4(W4TO22), .W5(W5TO22), .W6(W6TO22), .W7(W7TO22), .W8(W8TO22), .W9(W9TO22), .W10(W10TO22), .W11(W11TO22), .W12(W12TO22), .W13(W13TO22), .W14(W14TO22), .W15(W15TO22), .W16(W16TO22), .W17(W17TO22), .W18(W18TO22), .W19(W19TO22), .W20(W20TO22), .W21(W21TO22), .W22(W22TO22), .W23(W23TO22), .W24(W24TO22), .W25(W25TO22), .W26(W26TO22), .W27(W27TO22), .W28(W28TO22), .W29(W29TO22), .W30(W30TO22), .W31(W31TO22), .W32(W32TO22), .W33(W33TO22), .W34(W34TO22), .W35(W35TO22), .W36(W36TO22), .W37(W37TO22), .W38(W38TO22), .W39(W39TO22), .W40(W40TO22), .W41(W41TO22), .W42(W42TO22), .W43(W43TO22), .W44(W44TO22), .W45(W45TO22), .W46(W46TO22), .W47(W47TO22), .W48(W48TO22), .W49(W49TO22), .W50(W50TO22), .W51(W51TO22), .W52(W52TO22), .W53(W53TO22), .W54(W54TO22), .W55(W55TO22), .W56(W56TO22), .W57(W57TO22), .W58(W58TO22), .W59(W59TO22), .W60(W60TO22), .W61(W61TO22), .W62(W62TO22), .W63(W63TO22)) neuron22(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out22));
neuron64in #(.W0(W0TO23), .W1(W1TO23), .W2(W2TO23), .W3(W3TO23), .W4(W4TO23), .W5(W5TO23), .W6(W6TO23), .W7(W7TO23), .W8(W8TO23), .W9(W9TO23), .W10(W10TO23), .W11(W11TO23), .W12(W12TO23), .W13(W13TO23), .W14(W14TO23), .W15(W15TO23), .W16(W16TO23), .W17(W17TO23), .W18(W18TO23), .W19(W19TO23), .W20(W20TO23), .W21(W21TO23), .W22(W22TO23), .W23(W23TO23), .W24(W24TO23), .W25(W25TO23), .W26(W26TO23), .W27(W27TO23), .W28(W28TO23), .W29(W29TO23), .W30(W30TO23), .W31(W31TO23), .W32(W32TO23), .W33(W33TO23), .W34(W34TO23), .W35(W35TO23), .W36(W36TO23), .W37(W37TO23), .W38(W38TO23), .W39(W39TO23), .W40(W40TO23), .W41(W41TO23), .W42(W42TO23), .W43(W43TO23), .W44(W44TO23), .W45(W45TO23), .W46(W46TO23), .W47(W47TO23), .W48(W48TO23), .W49(W49TO23), .W50(W50TO23), .W51(W51TO23), .W52(W52TO23), .W53(W53TO23), .W54(W54TO23), .W55(W55TO23), .W56(W56TO23), .W57(W57TO23), .W58(W58TO23), .W59(W59TO23), .W60(W60TO23), .W61(W61TO23), .W62(W62TO23), .W63(W63TO23)) neuron23(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out23));
neuron64in #(.W0(W0TO24), .W1(W1TO24), .W2(W2TO24), .W3(W3TO24), .W4(W4TO24), .W5(W5TO24), .W6(W6TO24), .W7(W7TO24), .W8(W8TO24), .W9(W9TO24), .W10(W10TO24), .W11(W11TO24), .W12(W12TO24), .W13(W13TO24), .W14(W14TO24), .W15(W15TO24), .W16(W16TO24), .W17(W17TO24), .W18(W18TO24), .W19(W19TO24), .W20(W20TO24), .W21(W21TO24), .W22(W22TO24), .W23(W23TO24), .W24(W24TO24), .W25(W25TO24), .W26(W26TO24), .W27(W27TO24), .W28(W28TO24), .W29(W29TO24), .W30(W30TO24), .W31(W31TO24), .W32(W32TO24), .W33(W33TO24), .W34(W34TO24), .W35(W35TO24), .W36(W36TO24), .W37(W37TO24), .W38(W38TO24), .W39(W39TO24), .W40(W40TO24), .W41(W41TO24), .W42(W42TO24), .W43(W43TO24), .W44(W44TO24), .W45(W45TO24), .W46(W46TO24), .W47(W47TO24), .W48(W48TO24), .W49(W49TO24), .W50(W50TO24), .W51(W51TO24), .W52(W52TO24), .W53(W53TO24), .W54(W54TO24), .W55(W55TO24), .W56(W56TO24), .W57(W57TO24), .W58(W58TO24), .W59(W59TO24), .W60(W60TO24), .W61(W61TO24), .W62(W62TO24), .W63(W63TO24)) neuron24(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out24));
neuron64in #(.W0(W0TO25), .W1(W1TO25), .W2(W2TO25), .W3(W3TO25), .W4(W4TO25), .W5(W5TO25), .W6(W6TO25), .W7(W7TO25), .W8(W8TO25), .W9(W9TO25), .W10(W10TO25), .W11(W11TO25), .W12(W12TO25), .W13(W13TO25), .W14(W14TO25), .W15(W15TO25), .W16(W16TO25), .W17(W17TO25), .W18(W18TO25), .W19(W19TO25), .W20(W20TO25), .W21(W21TO25), .W22(W22TO25), .W23(W23TO25), .W24(W24TO25), .W25(W25TO25), .W26(W26TO25), .W27(W27TO25), .W28(W28TO25), .W29(W29TO25), .W30(W30TO25), .W31(W31TO25), .W32(W32TO25), .W33(W33TO25), .W34(W34TO25), .W35(W35TO25), .W36(W36TO25), .W37(W37TO25), .W38(W38TO25), .W39(W39TO25), .W40(W40TO25), .W41(W41TO25), .W42(W42TO25), .W43(W43TO25), .W44(W44TO25), .W45(W45TO25), .W46(W46TO25), .W47(W47TO25), .W48(W48TO25), .W49(W49TO25), .W50(W50TO25), .W51(W51TO25), .W52(W52TO25), .W53(W53TO25), .W54(W54TO25), .W55(W55TO25), .W56(W56TO25), .W57(W57TO25), .W58(W58TO25), .W59(W59TO25), .W60(W60TO25), .W61(W61TO25), .W62(W62TO25), .W63(W63TO25)) neuron25(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out25));
neuron64in #(.W0(W0TO26), .W1(W1TO26), .W2(W2TO26), .W3(W3TO26), .W4(W4TO26), .W5(W5TO26), .W6(W6TO26), .W7(W7TO26), .W8(W8TO26), .W9(W9TO26), .W10(W10TO26), .W11(W11TO26), .W12(W12TO26), .W13(W13TO26), .W14(W14TO26), .W15(W15TO26), .W16(W16TO26), .W17(W17TO26), .W18(W18TO26), .W19(W19TO26), .W20(W20TO26), .W21(W21TO26), .W22(W22TO26), .W23(W23TO26), .W24(W24TO26), .W25(W25TO26), .W26(W26TO26), .W27(W27TO26), .W28(W28TO26), .W29(W29TO26), .W30(W30TO26), .W31(W31TO26), .W32(W32TO26), .W33(W33TO26), .W34(W34TO26), .W35(W35TO26), .W36(W36TO26), .W37(W37TO26), .W38(W38TO26), .W39(W39TO26), .W40(W40TO26), .W41(W41TO26), .W42(W42TO26), .W43(W43TO26), .W44(W44TO26), .W45(W45TO26), .W46(W46TO26), .W47(W47TO26), .W48(W48TO26), .W49(W49TO26), .W50(W50TO26), .W51(W51TO26), .W52(W52TO26), .W53(W53TO26), .W54(W54TO26), .W55(W55TO26), .W56(W56TO26), .W57(W57TO26), .W58(W58TO26), .W59(W59TO26), .W60(W60TO26), .W61(W61TO26), .W62(W62TO26), .W63(W63TO26)) neuron26(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out26));
neuron64in #(.W0(W0TO27), .W1(W1TO27), .W2(W2TO27), .W3(W3TO27), .W4(W4TO27), .W5(W5TO27), .W6(W6TO27), .W7(W7TO27), .W8(W8TO27), .W9(W9TO27), .W10(W10TO27), .W11(W11TO27), .W12(W12TO27), .W13(W13TO27), .W14(W14TO27), .W15(W15TO27), .W16(W16TO27), .W17(W17TO27), .W18(W18TO27), .W19(W19TO27), .W20(W20TO27), .W21(W21TO27), .W22(W22TO27), .W23(W23TO27), .W24(W24TO27), .W25(W25TO27), .W26(W26TO27), .W27(W27TO27), .W28(W28TO27), .W29(W29TO27), .W30(W30TO27), .W31(W31TO27), .W32(W32TO27), .W33(W33TO27), .W34(W34TO27), .W35(W35TO27), .W36(W36TO27), .W37(W37TO27), .W38(W38TO27), .W39(W39TO27), .W40(W40TO27), .W41(W41TO27), .W42(W42TO27), .W43(W43TO27), .W44(W44TO27), .W45(W45TO27), .W46(W46TO27), .W47(W47TO27), .W48(W48TO27), .W49(W49TO27), .W50(W50TO27), .W51(W51TO27), .W52(W52TO27), .W53(W53TO27), .W54(W54TO27), .W55(W55TO27), .W56(W56TO27), .W57(W57TO27), .W58(W58TO27), .W59(W59TO27), .W60(W60TO27), .W61(W61TO27), .W62(W62TO27), .W63(W63TO27)) neuron27(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out27));
neuron64in #(.W0(W0TO28), .W1(W1TO28), .W2(W2TO28), .W3(W3TO28), .W4(W4TO28), .W5(W5TO28), .W6(W6TO28), .W7(W7TO28), .W8(W8TO28), .W9(W9TO28), .W10(W10TO28), .W11(W11TO28), .W12(W12TO28), .W13(W13TO28), .W14(W14TO28), .W15(W15TO28), .W16(W16TO28), .W17(W17TO28), .W18(W18TO28), .W19(W19TO28), .W20(W20TO28), .W21(W21TO28), .W22(W22TO28), .W23(W23TO28), .W24(W24TO28), .W25(W25TO28), .W26(W26TO28), .W27(W27TO28), .W28(W28TO28), .W29(W29TO28), .W30(W30TO28), .W31(W31TO28), .W32(W32TO28), .W33(W33TO28), .W34(W34TO28), .W35(W35TO28), .W36(W36TO28), .W37(W37TO28), .W38(W38TO28), .W39(W39TO28), .W40(W40TO28), .W41(W41TO28), .W42(W42TO28), .W43(W43TO28), .W44(W44TO28), .W45(W45TO28), .W46(W46TO28), .W47(W47TO28), .W48(W48TO28), .W49(W49TO28), .W50(W50TO28), .W51(W51TO28), .W52(W52TO28), .W53(W53TO28), .W54(W54TO28), .W55(W55TO28), .W56(W56TO28), .W57(W57TO28), .W58(W58TO28), .W59(W59TO28), .W60(W60TO28), .W61(W61TO28), .W62(W62TO28), .W63(W63TO28)) neuron28(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out28));
neuron64in #(.W0(W0TO29), .W1(W1TO29), .W2(W2TO29), .W3(W3TO29), .W4(W4TO29), .W5(W5TO29), .W6(W6TO29), .W7(W7TO29), .W8(W8TO29), .W9(W9TO29), .W10(W10TO29), .W11(W11TO29), .W12(W12TO29), .W13(W13TO29), .W14(W14TO29), .W15(W15TO29), .W16(W16TO29), .W17(W17TO29), .W18(W18TO29), .W19(W19TO29), .W20(W20TO29), .W21(W21TO29), .W22(W22TO29), .W23(W23TO29), .W24(W24TO29), .W25(W25TO29), .W26(W26TO29), .W27(W27TO29), .W28(W28TO29), .W29(W29TO29), .W30(W30TO29), .W31(W31TO29), .W32(W32TO29), .W33(W33TO29), .W34(W34TO29), .W35(W35TO29), .W36(W36TO29), .W37(W37TO29), .W38(W38TO29), .W39(W39TO29), .W40(W40TO29), .W41(W41TO29), .W42(W42TO29), .W43(W43TO29), .W44(W44TO29), .W45(W45TO29), .W46(W46TO29), .W47(W47TO29), .W48(W48TO29), .W49(W49TO29), .W50(W50TO29), .W51(W51TO29), .W52(W52TO29), .W53(W53TO29), .W54(W54TO29), .W55(W55TO29), .W56(W56TO29), .W57(W57TO29), .W58(W58TO29), .W59(W59TO29), .W60(W60TO29), .W61(W61TO29), .W62(W62TO29), .W63(W63TO29)) neuron29(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out29));
neuron64in #(.W0(W0TO30), .W1(W1TO30), .W2(W2TO30), .W3(W3TO30), .W4(W4TO30), .W5(W5TO30), .W6(W6TO30), .W7(W7TO30), .W8(W8TO30), .W9(W9TO30), .W10(W10TO30), .W11(W11TO30), .W12(W12TO30), .W13(W13TO30), .W14(W14TO30), .W15(W15TO30), .W16(W16TO30), .W17(W17TO30), .W18(W18TO30), .W19(W19TO30), .W20(W20TO30), .W21(W21TO30), .W22(W22TO30), .W23(W23TO30), .W24(W24TO30), .W25(W25TO30), .W26(W26TO30), .W27(W27TO30), .W28(W28TO30), .W29(W29TO30), .W30(W30TO30), .W31(W31TO30), .W32(W32TO30), .W33(W33TO30), .W34(W34TO30), .W35(W35TO30), .W36(W36TO30), .W37(W37TO30), .W38(W38TO30), .W39(W39TO30), .W40(W40TO30), .W41(W41TO30), .W42(W42TO30), .W43(W43TO30), .W44(W44TO30), .W45(W45TO30), .W46(W46TO30), .W47(W47TO30), .W48(W48TO30), .W49(W49TO30), .W50(W50TO30), .W51(W51TO30), .W52(W52TO30), .W53(W53TO30), .W54(W54TO30), .W55(W55TO30), .W56(W56TO30), .W57(W57TO30), .W58(W58TO30), .W59(W59TO30), .W60(W60TO30), .W61(W61TO30), .W62(W62TO30), .W63(W63TO30)) neuron30(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out30));
neuron64in #(.W0(W0TO31), .W1(W1TO31), .W2(W2TO31), .W3(W3TO31), .W4(W4TO31), .W5(W5TO31), .W6(W6TO31), .W7(W7TO31), .W8(W8TO31), .W9(W9TO31), .W10(W10TO31), .W11(W11TO31), .W12(W12TO31), .W13(W13TO31), .W14(W14TO31), .W15(W15TO31), .W16(W16TO31), .W17(W17TO31), .W18(W18TO31), .W19(W19TO31), .W20(W20TO31), .W21(W21TO31), .W22(W22TO31), .W23(W23TO31), .W24(W24TO31), .W25(W25TO31), .W26(W26TO31), .W27(W27TO31), .W28(W28TO31), .W29(W29TO31), .W30(W30TO31), .W31(W31TO31), .W32(W32TO31), .W33(W33TO31), .W34(W34TO31), .W35(W35TO31), .W36(W36TO31), .W37(W37TO31), .W38(W38TO31), .W39(W39TO31), .W40(W40TO31), .W41(W41TO31), .W42(W42TO31), .W43(W43TO31), .W44(W44TO31), .W45(W45TO31), .W46(W46TO31), .W47(W47TO31), .W48(W48TO31), .W49(W49TO31), .W50(W50TO31), .W51(W51TO31), .W52(W52TO31), .W53(W53TO31), .W54(W54TO31), .W55(W55TO31), .W56(W56TO31), .W57(W57TO31), .W58(W58TO31), .W59(W59TO31), .W60(W60TO31), .W61(W61TO31), .W62(W62TO31), .W63(W63TO31)) neuron31(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out31));
neuron64in #(.W0(W0TO32), .W1(W1TO32), .W2(W2TO32), .W3(W3TO32), .W4(W4TO32), .W5(W5TO32), .W6(W6TO32), .W7(W7TO32), .W8(W8TO32), .W9(W9TO32), .W10(W10TO32), .W11(W11TO32), .W12(W12TO32), .W13(W13TO32), .W14(W14TO32), .W15(W15TO32), .W16(W16TO32), .W17(W17TO32), .W18(W18TO32), .W19(W19TO32), .W20(W20TO32), .W21(W21TO32), .W22(W22TO32), .W23(W23TO32), .W24(W24TO32), .W25(W25TO32), .W26(W26TO32), .W27(W27TO32), .W28(W28TO32), .W29(W29TO32), .W30(W30TO32), .W31(W31TO32), .W32(W32TO32), .W33(W33TO32), .W34(W34TO32), .W35(W35TO32), .W36(W36TO32), .W37(W37TO32), .W38(W38TO32), .W39(W39TO32), .W40(W40TO32), .W41(W41TO32), .W42(W42TO32), .W43(W43TO32), .W44(W44TO32), .W45(W45TO32), .W46(W46TO32), .W47(W47TO32), .W48(W48TO32), .W49(W49TO32), .W50(W50TO32), .W51(W51TO32), .W52(W52TO32), .W53(W53TO32), .W54(W54TO32), .W55(W55TO32), .W56(W56TO32), .W57(W57TO32), .W58(W58TO32), .W59(W59TO32), .W60(W60TO32), .W61(W61TO32), .W62(W62TO32), .W63(W63TO32)) neuron32(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out32));
neuron64in #(.W0(W0TO33), .W1(W1TO33), .W2(W2TO33), .W3(W3TO33), .W4(W4TO33), .W5(W5TO33), .W6(W6TO33), .W7(W7TO33), .W8(W8TO33), .W9(W9TO33), .W10(W10TO33), .W11(W11TO33), .W12(W12TO33), .W13(W13TO33), .W14(W14TO33), .W15(W15TO33), .W16(W16TO33), .W17(W17TO33), .W18(W18TO33), .W19(W19TO33), .W20(W20TO33), .W21(W21TO33), .W22(W22TO33), .W23(W23TO33), .W24(W24TO33), .W25(W25TO33), .W26(W26TO33), .W27(W27TO33), .W28(W28TO33), .W29(W29TO33), .W30(W30TO33), .W31(W31TO33), .W32(W32TO33), .W33(W33TO33), .W34(W34TO33), .W35(W35TO33), .W36(W36TO33), .W37(W37TO33), .W38(W38TO33), .W39(W39TO33), .W40(W40TO33), .W41(W41TO33), .W42(W42TO33), .W43(W43TO33), .W44(W44TO33), .W45(W45TO33), .W46(W46TO33), .W47(W47TO33), .W48(W48TO33), .W49(W49TO33), .W50(W50TO33), .W51(W51TO33), .W52(W52TO33), .W53(W53TO33), .W54(W54TO33), .W55(W55TO33), .W56(W56TO33), .W57(W57TO33), .W58(W58TO33), .W59(W59TO33), .W60(W60TO33), .W61(W61TO33), .W62(W62TO33), .W63(W63TO33)) neuron33(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out33));
neuron64in #(.W0(W0TO34), .W1(W1TO34), .W2(W2TO34), .W3(W3TO34), .W4(W4TO34), .W5(W5TO34), .W6(W6TO34), .W7(W7TO34), .W8(W8TO34), .W9(W9TO34), .W10(W10TO34), .W11(W11TO34), .W12(W12TO34), .W13(W13TO34), .W14(W14TO34), .W15(W15TO34), .W16(W16TO34), .W17(W17TO34), .W18(W18TO34), .W19(W19TO34), .W20(W20TO34), .W21(W21TO34), .W22(W22TO34), .W23(W23TO34), .W24(W24TO34), .W25(W25TO34), .W26(W26TO34), .W27(W27TO34), .W28(W28TO34), .W29(W29TO34), .W30(W30TO34), .W31(W31TO34), .W32(W32TO34), .W33(W33TO34), .W34(W34TO34), .W35(W35TO34), .W36(W36TO34), .W37(W37TO34), .W38(W38TO34), .W39(W39TO34), .W40(W40TO34), .W41(W41TO34), .W42(W42TO34), .W43(W43TO34), .W44(W44TO34), .W45(W45TO34), .W46(W46TO34), .W47(W47TO34), .W48(W48TO34), .W49(W49TO34), .W50(W50TO34), .W51(W51TO34), .W52(W52TO34), .W53(W53TO34), .W54(W54TO34), .W55(W55TO34), .W56(W56TO34), .W57(W57TO34), .W58(W58TO34), .W59(W59TO34), .W60(W60TO34), .W61(W61TO34), .W62(W62TO34), .W63(W63TO34)) neuron34(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out34));
neuron64in #(.W0(W0TO35), .W1(W1TO35), .W2(W2TO35), .W3(W3TO35), .W4(W4TO35), .W5(W5TO35), .W6(W6TO35), .W7(W7TO35), .W8(W8TO35), .W9(W9TO35), .W10(W10TO35), .W11(W11TO35), .W12(W12TO35), .W13(W13TO35), .W14(W14TO35), .W15(W15TO35), .W16(W16TO35), .W17(W17TO35), .W18(W18TO35), .W19(W19TO35), .W20(W20TO35), .W21(W21TO35), .W22(W22TO35), .W23(W23TO35), .W24(W24TO35), .W25(W25TO35), .W26(W26TO35), .W27(W27TO35), .W28(W28TO35), .W29(W29TO35), .W30(W30TO35), .W31(W31TO35), .W32(W32TO35), .W33(W33TO35), .W34(W34TO35), .W35(W35TO35), .W36(W36TO35), .W37(W37TO35), .W38(W38TO35), .W39(W39TO35), .W40(W40TO35), .W41(W41TO35), .W42(W42TO35), .W43(W43TO35), .W44(W44TO35), .W45(W45TO35), .W46(W46TO35), .W47(W47TO35), .W48(W48TO35), .W49(W49TO35), .W50(W50TO35), .W51(W51TO35), .W52(W52TO35), .W53(W53TO35), .W54(W54TO35), .W55(W55TO35), .W56(W56TO35), .W57(W57TO35), .W58(W58TO35), .W59(W59TO35), .W60(W60TO35), .W61(W61TO35), .W62(W62TO35), .W63(W63TO35)) neuron35(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out35));
neuron64in #(.W0(W0TO36), .W1(W1TO36), .W2(W2TO36), .W3(W3TO36), .W4(W4TO36), .W5(W5TO36), .W6(W6TO36), .W7(W7TO36), .W8(W8TO36), .W9(W9TO36), .W10(W10TO36), .W11(W11TO36), .W12(W12TO36), .W13(W13TO36), .W14(W14TO36), .W15(W15TO36), .W16(W16TO36), .W17(W17TO36), .W18(W18TO36), .W19(W19TO36), .W20(W20TO36), .W21(W21TO36), .W22(W22TO36), .W23(W23TO36), .W24(W24TO36), .W25(W25TO36), .W26(W26TO36), .W27(W27TO36), .W28(W28TO36), .W29(W29TO36), .W30(W30TO36), .W31(W31TO36), .W32(W32TO36), .W33(W33TO36), .W34(W34TO36), .W35(W35TO36), .W36(W36TO36), .W37(W37TO36), .W38(W38TO36), .W39(W39TO36), .W40(W40TO36), .W41(W41TO36), .W42(W42TO36), .W43(W43TO36), .W44(W44TO36), .W45(W45TO36), .W46(W46TO36), .W47(W47TO36), .W48(W48TO36), .W49(W49TO36), .W50(W50TO36), .W51(W51TO36), .W52(W52TO36), .W53(W53TO36), .W54(W54TO36), .W55(W55TO36), .W56(W56TO36), .W57(W57TO36), .W58(W58TO36), .W59(W59TO36), .W60(W60TO36), .W61(W61TO36), .W62(W62TO36), .W63(W63TO36)) neuron36(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out36));
neuron64in #(.W0(W0TO37), .W1(W1TO37), .W2(W2TO37), .W3(W3TO37), .W4(W4TO37), .W5(W5TO37), .W6(W6TO37), .W7(W7TO37), .W8(W8TO37), .W9(W9TO37), .W10(W10TO37), .W11(W11TO37), .W12(W12TO37), .W13(W13TO37), .W14(W14TO37), .W15(W15TO37), .W16(W16TO37), .W17(W17TO37), .W18(W18TO37), .W19(W19TO37), .W20(W20TO37), .W21(W21TO37), .W22(W22TO37), .W23(W23TO37), .W24(W24TO37), .W25(W25TO37), .W26(W26TO37), .W27(W27TO37), .W28(W28TO37), .W29(W29TO37), .W30(W30TO37), .W31(W31TO37), .W32(W32TO37), .W33(W33TO37), .W34(W34TO37), .W35(W35TO37), .W36(W36TO37), .W37(W37TO37), .W38(W38TO37), .W39(W39TO37), .W40(W40TO37), .W41(W41TO37), .W42(W42TO37), .W43(W43TO37), .W44(W44TO37), .W45(W45TO37), .W46(W46TO37), .W47(W47TO37), .W48(W48TO37), .W49(W49TO37), .W50(W50TO37), .W51(W51TO37), .W52(W52TO37), .W53(W53TO37), .W54(W54TO37), .W55(W55TO37), .W56(W56TO37), .W57(W57TO37), .W58(W58TO37), .W59(W59TO37), .W60(W60TO37), .W61(W61TO37), .W62(W62TO37), .W63(W63TO37)) neuron37(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out37));
neuron64in #(.W0(W0TO38), .W1(W1TO38), .W2(W2TO38), .W3(W3TO38), .W4(W4TO38), .W5(W5TO38), .W6(W6TO38), .W7(W7TO38), .W8(W8TO38), .W9(W9TO38), .W10(W10TO38), .W11(W11TO38), .W12(W12TO38), .W13(W13TO38), .W14(W14TO38), .W15(W15TO38), .W16(W16TO38), .W17(W17TO38), .W18(W18TO38), .W19(W19TO38), .W20(W20TO38), .W21(W21TO38), .W22(W22TO38), .W23(W23TO38), .W24(W24TO38), .W25(W25TO38), .W26(W26TO38), .W27(W27TO38), .W28(W28TO38), .W29(W29TO38), .W30(W30TO38), .W31(W31TO38), .W32(W32TO38), .W33(W33TO38), .W34(W34TO38), .W35(W35TO38), .W36(W36TO38), .W37(W37TO38), .W38(W38TO38), .W39(W39TO38), .W40(W40TO38), .W41(W41TO38), .W42(W42TO38), .W43(W43TO38), .W44(W44TO38), .W45(W45TO38), .W46(W46TO38), .W47(W47TO38), .W48(W48TO38), .W49(W49TO38), .W50(W50TO38), .W51(W51TO38), .W52(W52TO38), .W53(W53TO38), .W54(W54TO38), .W55(W55TO38), .W56(W56TO38), .W57(W57TO38), .W58(W58TO38), .W59(W59TO38), .W60(W60TO38), .W61(W61TO38), .W62(W62TO38), .W63(W63TO38)) neuron38(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out38));
neuron64in #(.W0(W0TO39), .W1(W1TO39), .W2(W2TO39), .W3(W3TO39), .W4(W4TO39), .W5(W5TO39), .W6(W6TO39), .W7(W7TO39), .W8(W8TO39), .W9(W9TO39), .W10(W10TO39), .W11(W11TO39), .W12(W12TO39), .W13(W13TO39), .W14(W14TO39), .W15(W15TO39), .W16(W16TO39), .W17(W17TO39), .W18(W18TO39), .W19(W19TO39), .W20(W20TO39), .W21(W21TO39), .W22(W22TO39), .W23(W23TO39), .W24(W24TO39), .W25(W25TO39), .W26(W26TO39), .W27(W27TO39), .W28(W28TO39), .W29(W29TO39), .W30(W30TO39), .W31(W31TO39), .W32(W32TO39), .W33(W33TO39), .W34(W34TO39), .W35(W35TO39), .W36(W36TO39), .W37(W37TO39), .W38(W38TO39), .W39(W39TO39), .W40(W40TO39), .W41(W41TO39), .W42(W42TO39), .W43(W43TO39), .W44(W44TO39), .W45(W45TO39), .W46(W46TO39), .W47(W47TO39), .W48(W48TO39), .W49(W49TO39), .W50(W50TO39), .W51(W51TO39), .W52(W52TO39), .W53(W53TO39), .W54(W54TO39), .W55(W55TO39), .W56(W56TO39), .W57(W57TO39), .W58(W58TO39), .W59(W59TO39), .W60(W60TO39), .W61(W61TO39), .W62(W62TO39), .W63(W63TO39)) neuron39(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out39));
neuron64in #(.W0(W0TO40), .W1(W1TO40), .W2(W2TO40), .W3(W3TO40), .W4(W4TO40), .W5(W5TO40), .W6(W6TO40), .W7(W7TO40), .W8(W8TO40), .W9(W9TO40), .W10(W10TO40), .W11(W11TO40), .W12(W12TO40), .W13(W13TO40), .W14(W14TO40), .W15(W15TO40), .W16(W16TO40), .W17(W17TO40), .W18(W18TO40), .W19(W19TO40), .W20(W20TO40), .W21(W21TO40), .W22(W22TO40), .W23(W23TO40), .W24(W24TO40), .W25(W25TO40), .W26(W26TO40), .W27(W27TO40), .W28(W28TO40), .W29(W29TO40), .W30(W30TO40), .W31(W31TO40), .W32(W32TO40), .W33(W33TO40), .W34(W34TO40), .W35(W35TO40), .W36(W36TO40), .W37(W37TO40), .W38(W38TO40), .W39(W39TO40), .W40(W40TO40), .W41(W41TO40), .W42(W42TO40), .W43(W43TO40), .W44(W44TO40), .W45(W45TO40), .W46(W46TO40), .W47(W47TO40), .W48(W48TO40), .W49(W49TO40), .W50(W50TO40), .W51(W51TO40), .W52(W52TO40), .W53(W53TO40), .W54(W54TO40), .W55(W55TO40), .W56(W56TO40), .W57(W57TO40), .W58(W58TO40), .W59(W59TO40), .W60(W60TO40), .W61(W61TO40), .W62(W62TO40), .W63(W63TO40)) neuron40(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out40));
neuron64in #(.W0(W0TO41), .W1(W1TO41), .W2(W2TO41), .W3(W3TO41), .W4(W4TO41), .W5(W5TO41), .W6(W6TO41), .W7(W7TO41), .W8(W8TO41), .W9(W9TO41), .W10(W10TO41), .W11(W11TO41), .W12(W12TO41), .W13(W13TO41), .W14(W14TO41), .W15(W15TO41), .W16(W16TO41), .W17(W17TO41), .W18(W18TO41), .W19(W19TO41), .W20(W20TO41), .W21(W21TO41), .W22(W22TO41), .W23(W23TO41), .W24(W24TO41), .W25(W25TO41), .W26(W26TO41), .W27(W27TO41), .W28(W28TO41), .W29(W29TO41), .W30(W30TO41), .W31(W31TO41), .W32(W32TO41), .W33(W33TO41), .W34(W34TO41), .W35(W35TO41), .W36(W36TO41), .W37(W37TO41), .W38(W38TO41), .W39(W39TO41), .W40(W40TO41), .W41(W41TO41), .W42(W42TO41), .W43(W43TO41), .W44(W44TO41), .W45(W45TO41), .W46(W46TO41), .W47(W47TO41), .W48(W48TO41), .W49(W49TO41), .W50(W50TO41), .W51(W51TO41), .W52(W52TO41), .W53(W53TO41), .W54(W54TO41), .W55(W55TO41), .W56(W56TO41), .W57(W57TO41), .W58(W58TO41), .W59(W59TO41), .W60(W60TO41), .W61(W61TO41), .W62(W62TO41), .W63(W63TO41)) neuron41(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out41));
neuron64in #(.W0(W0TO42), .W1(W1TO42), .W2(W2TO42), .W3(W3TO42), .W4(W4TO42), .W5(W5TO42), .W6(W6TO42), .W7(W7TO42), .W8(W8TO42), .W9(W9TO42), .W10(W10TO42), .W11(W11TO42), .W12(W12TO42), .W13(W13TO42), .W14(W14TO42), .W15(W15TO42), .W16(W16TO42), .W17(W17TO42), .W18(W18TO42), .W19(W19TO42), .W20(W20TO42), .W21(W21TO42), .W22(W22TO42), .W23(W23TO42), .W24(W24TO42), .W25(W25TO42), .W26(W26TO42), .W27(W27TO42), .W28(W28TO42), .W29(W29TO42), .W30(W30TO42), .W31(W31TO42), .W32(W32TO42), .W33(W33TO42), .W34(W34TO42), .W35(W35TO42), .W36(W36TO42), .W37(W37TO42), .W38(W38TO42), .W39(W39TO42), .W40(W40TO42), .W41(W41TO42), .W42(W42TO42), .W43(W43TO42), .W44(W44TO42), .W45(W45TO42), .W46(W46TO42), .W47(W47TO42), .W48(W48TO42), .W49(W49TO42), .W50(W50TO42), .W51(W51TO42), .W52(W52TO42), .W53(W53TO42), .W54(W54TO42), .W55(W55TO42), .W56(W56TO42), .W57(W57TO42), .W58(W58TO42), .W59(W59TO42), .W60(W60TO42), .W61(W61TO42), .W62(W62TO42), .W63(W63TO42)) neuron42(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out42));
neuron64in #(.W0(W0TO43), .W1(W1TO43), .W2(W2TO43), .W3(W3TO43), .W4(W4TO43), .W5(W5TO43), .W6(W6TO43), .W7(W7TO43), .W8(W8TO43), .W9(W9TO43), .W10(W10TO43), .W11(W11TO43), .W12(W12TO43), .W13(W13TO43), .W14(W14TO43), .W15(W15TO43), .W16(W16TO43), .W17(W17TO43), .W18(W18TO43), .W19(W19TO43), .W20(W20TO43), .W21(W21TO43), .W22(W22TO43), .W23(W23TO43), .W24(W24TO43), .W25(W25TO43), .W26(W26TO43), .W27(W27TO43), .W28(W28TO43), .W29(W29TO43), .W30(W30TO43), .W31(W31TO43), .W32(W32TO43), .W33(W33TO43), .W34(W34TO43), .W35(W35TO43), .W36(W36TO43), .W37(W37TO43), .W38(W38TO43), .W39(W39TO43), .W40(W40TO43), .W41(W41TO43), .W42(W42TO43), .W43(W43TO43), .W44(W44TO43), .W45(W45TO43), .W46(W46TO43), .W47(W47TO43), .W48(W48TO43), .W49(W49TO43), .W50(W50TO43), .W51(W51TO43), .W52(W52TO43), .W53(W53TO43), .W54(W54TO43), .W55(W55TO43), .W56(W56TO43), .W57(W57TO43), .W58(W58TO43), .W59(W59TO43), .W60(W60TO43), .W61(W61TO43), .W62(W62TO43), .W63(W63TO43)) neuron43(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out43));
neuron64in #(.W0(W0TO44), .W1(W1TO44), .W2(W2TO44), .W3(W3TO44), .W4(W4TO44), .W5(W5TO44), .W6(W6TO44), .W7(W7TO44), .W8(W8TO44), .W9(W9TO44), .W10(W10TO44), .W11(W11TO44), .W12(W12TO44), .W13(W13TO44), .W14(W14TO44), .W15(W15TO44), .W16(W16TO44), .W17(W17TO44), .W18(W18TO44), .W19(W19TO44), .W20(W20TO44), .W21(W21TO44), .W22(W22TO44), .W23(W23TO44), .W24(W24TO44), .W25(W25TO44), .W26(W26TO44), .W27(W27TO44), .W28(W28TO44), .W29(W29TO44), .W30(W30TO44), .W31(W31TO44), .W32(W32TO44), .W33(W33TO44), .W34(W34TO44), .W35(W35TO44), .W36(W36TO44), .W37(W37TO44), .W38(W38TO44), .W39(W39TO44), .W40(W40TO44), .W41(W41TO44), .W42(W42TO44), .W43(W43TO44), .W44(W44TO44), .W45(W45TO44), .W46(W46TO44), .W47(W47TO44), .W48(W48TO44), .W49(W49TO44), .W50(W50TO44), .W51(W51TO44), .W52(W52TO44), .W53(W53TO44), .W54(W54TO44), .W55(W55TO44), .W56(W56TO44), .W57(W57TO44), .W58(W58TO44), .W59(W59TO44), .W60(W60TO44), .W61(W61TO44), .W62(W62TO44), .W63(W63TO44)) neuron44(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out44));
neuron64in #(.W0(W0TO45), .W1(W1TO45), .W2(W2TO45), .W3(W3TO45), .W4(W4TO45), .W5(W5TO45), .W6(W6TO45), .W7(W7TO45), .W8(W8TO45), .W9(W9TO45), .W10(W10TO45), .W11(W11TO45), .W12(W12TO45), .W13(W13TO45), .W14(W14TO45), .W15(W15TO45), .W16(W16TO45), .W17(W17TO45), .W18(W18TO45), .W19(W19TO45), .W20(W20TO45), .W21(W21TO45), .W22(W22TO45), .W23(W23TO45), .W24(W24TO45), .W25(W25TO45), .W26(W26TO45), .W27(W27TO45), .W28(W28TO45), .W29(W29TO45), .W30(W30TO45), .W31(W31TO45), .W32(W32TO45), .W33(W33TO45), .W34(W34TO45), .W35(W35TO45), .W36(W36TO45), .W37(W37TO45), .W38(W38TO45), .W39(W39TO45), .W40(W40TO45), .W41(W41TO45), .W42(W42TO45), .W43(W43TO45), .W44(W44TO45), .W45(W45TO45), .W46(W46TO45), .W47(W47TO45), .W48(W48TO45), .W49(W49TO45), .W50(W50TO45), .W51(W51TO45), .W52(W52TO45), .W53(W53TO45), .W54(W54TO45), .W55(W55TO45), .W56(W56TO45), .W57(W57TO45), .W58(W58TO45), .W59(W59TO45), .W60(W60TO45), .W61(W61TO45), .W62(W62TO45), .W63(W63TO45)) neuron45(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out45));
neuron64in #(.W0(W0TO46), .W1(W1TO46), .W2(W2TO46), .W3(W3TO46), .W4(W4TO46), .W5(W5TO46), .W6(W6TO46), .W7(W7TO46), .W8(W8TO46), .W9(W9TO46), .W10(W10TO46), .W11(W11TO46), .W12(W12TO46), .W13(W13TO46), .W14(W14TO46), .W15(W15TO46), .W16(W16TO46), .W17(W17TO46), .W18(W18TO46), .W19(W19TO46), .W20(W20TO46), .W21(W21TO46), .W22(W22TO46), .W23(W23TO46), .W24(W24TO46), .W25(W25TO46), .W26(W26TO46), .W27(W27TO46), .W28(W28TO46), .W29(W29TO46), .W30(W30TO46), .W31(W31TO46), .W32(W32TO46), .W33(W33TO46), .W34(W34TO46), .W35(W35TO46), .W36(W36TO46), .W37(W37TO46), .W38(W38TO46), .W39(W39TO46), .W40(W40TO46), .W41(W41TO46), .W42(W42TO46), .W43(W43TO46), .W44(W44TO46), .W45(W45TO46), .W46(W46TO46), .W47(W47TO46), .W48(W48TO46), .W49(W49TO46), .W50(W50TO46), .W51(W51TO46), .W52(W52TO46), .W53(W53TO46), .W54(W54TO46), .W55(W55TO46), .W56(W56TO46), .W57(W57TO46), .W58(W58TO46), .W59(W59TO46), .W60(W60TO46), .W61(W61TO46), .W62(W62TO46), .W63(W63TO46)) neuron46(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out46));
neuron64in #(.W0(W0TO47), .W1(W1TO47), .W2(W2TO47), .W3(W3TO47), .W4(W4TO47), .W5(W5TO47), .W6(W6TO47), .W7(W7TO47), .W8(W8TO47), .W9(W9TO47), .W10(W10TO47), .W11(W11TO47), .W12(W12TO47), .W13(W13TO47), .W14(W14TO47), .W15(W15TO47), .W16(W16TO47), .W17(W17TO47), .W18(W18TO47), .W19(W19TO47), .W20(W20TO47), .W21(W21TO47), .W22(W22TO47), .W23(W23TO47), .W24(W24TO47), .W25(W25TO47), .W26(W26TO47), .W27(W27TO47), .W28(W28TO47), .W29(W29TO47), .W30(W30TO47), .W31(W31TO47), .W32(W32TO47), .W33(W33TO47), .W34(W34TO47), .W35(W35TO47), .W36(W36TO47), .W37(W37TO47), .W38(W38TO47), .W39(W39TO47), .W40(W40TO47), .W41(W41TO47), .W42(W42TO47), .W43(W43TO47), .W44(W44TO47), .W45(W45TO47), .W46(W46TO47), .W47(W47TO47), .W48(W48TO47), .W49(W49TO47), .W50(W50TO47), .W51(W51TO47), .W52(W52TO47), .W53(W53TO47), .W54(W54TO47), .W55(W55TO47), .W56(W56TO47), .W57(W57TO47), .W58(W58TO47), .W59(W59TO47), .W60(W60TO47), .W61(W61TO47), .W62(W62TO47), .W63(W63TO47)) neuron47(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out47));
neuron64in #(.W0(W0TO48), .W1(W1TO48), .W2(W2TO48), .W3(W3TO48), .W4(W4TO48), .W5(W5TO48), .W6(W6TO48), .W7(W7TO48), .W8(W8TO48), .W9(W9TO48), .W10(W10TO48), .W11(W11TO48), .W12(W12TO48), .W13(W13TO48), .W14(W14TO48), .W15(W15TO48), .W16(W16TO48), .W17(W17TO48), .W18(W18TO48), .W19(W19TO48), .W20(W20TO48), .W21(W21TO48), .W22(W22TO48), .W23(W23TO48), .W24(W24TO48), .W25(W25TO48), .W26(W26TO48), .W27(W27TO48), .W28(W28TO48), .W29(W29TO48), .W30(W30TO48), .W31(W31TO48), .W32(W32TO48), .W33(W33TO48), .W34(W34TO48), .W35(W35TO48), .W36(W36TO48), .W37(W37TO48), .W38(W38TO48), .W39(W39TO48), .W40(W40TO48), .W41(W41TO48), .W42(W42TO48), .W43(W43TO48), .W44(W44TO48), .W45(W45TO48), .W46(W46TO48), .W47(W47TO48), .W48(W48TO48), .W49(W49TO48), .W50(W50TO48), .W51(W51TO48), .W52(W52TO48), .W53(W53TO48), .W54(W54TO48), .W55(W55TO48), .W56(W56TO48), .W57(W57TO48), .W58(W58TO48), .W59(W59TO48), .W60(W60TO48), .W61(W61TO48), .W62(W62TO48), .W63(W63TO48)) neuron48(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out48));
neuron64in #(.W0(W0TO49), .W1(W1TO49), .W2(W2TO49), .W3(W3TO49), .W4(W4TO49), .W5(W5TO49), .W6(W6TO49), .W7(W7TO49), .W8(W8TO49), .W9(W9TO49), .W10(W10TO49), .W11(W11TO49), .W12(W12TO49), .W13(W13TO49), .W14(W14TO49), .W15(W15TO49), .W16(W16TO49), .W17(W17TO49), .W18(W18TO49), .W19(W19TO49), .W20(W20TO49), .W21(W21TO49), .W22(W22TO49), .W23(W23TO49), .W24(W24TO49), .W25(W25TO49), .W26(W26TO49), .W27(W27TO49), .W28(W28TO49), .W29(W29TO49), .W30(W30TO49), .W31(W31TO49), .W32(W32TO49), .W33(W33TO49), .W34(W34TO49), .W35(W35TO49), .W36(W36TO49), .W37(W37TO49), .W38(W38TO49), .W39(W39TO49), .W40(W40TO49), .W41(W41TO49), .W42(W42TO49), .W43(W43TO49), .W44(W44TO49), .W45(W45TO49), .W46(W46TO49), .W47(W47TO49), .W48(W48TO49), .W49(W49TO49), .W50(W50TO49), .W51(W51TO49), .W52(W52TO49), .W53(W53TO49), .W54(W54TO49), .W55(W55TO49), .W56(W56TO49), .W57(W57TO49), .W58(W58TO49), .W59(W59TO49), .W60(W60TO49), .W61(W61TO49), .W62(W62TO49), .W63(W63TO49)) neuron49(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out49));
neuron64in #(.W0(W0TO50), .W1(W1TO50), .W2(W2TO50), .W3(W3TO50), .W4(W4TO50), .W5(W5TO50), .W6(W6TO50), .W7(W7TO50), .W8(W8TO50), .W9(W9TO50), .W10(W10TO50), .W11(W11TO50), .W12(W12TO50), .W13(W13TO50), .W14(W14TO50), .W15(W15TO50), .W16(W16TO50), .W17(W17TO50), .W18(W18TO50), .W19(W19TO50), .W20(W20TO50), .W21(W21TO50), .W22(W22TO50), .W23(W23TO50), .W24(W24TO50), .W25(W25TO50), .W26(W26TO50), .W27(W27TO50), .W28(W28TO50), .W29(W29TO50), .W30(W30TO50), .W31(W31TO50), .W32(W32TO50), .W33(W33TO50), .W34(W34TO50), .W35(W35TO50), .W36(W36TO50), .W37(W37TO50), .W38(W38TO50), .W39(W39TO50), .W40(W40TO50), .W41(W41TO50), .W42(W42TO50), .W43(W43TO50), .W44(W44TO50), .W45(W45TO50), .W46(W46TO50), .W47(W47TO50), .W48(W48TO50), .W49(W49TO50), .W50(W50TO50), .W51(W51TO50), .W52(W52TO50), .W53(W53TO50), .W54(W54TO50), .W55(W55TO50), .W56(W56TO50), .W57(W57TO50), .W58(W58TO50), .W59(W59TO50), .W60(W60TO50), .W61(W61TO50), .W62(W62TO50), .W63(W63TO50)) neuron50(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out50));
neuron64in #(.W0(W0TO51), .W1(W1TO51), .W2(W2TO51), .W3(W3TO51), .W4(W4TO51), .W5(W5TO51), .W6(W6TO51), .W7(W7TO51), .W8(W8TO51), .W9(W9TO51), .W10(W10TO51), .W11(W11TO51), .W12(W12TO51), .W13(W13TO51), .W14(W14TO51), .W15(W15TO51), .W16(W16TO51), .W17(W17TO51), .W18(W18TO51), .W19(W19TO51), .W20(W20TO51), .W21(W21TO51), .W22(W22TO51), .W23(W23TO51), .W24(W24TO51), .W25(W25TO51), .W26(W26TO51), .W27(W27TO51), .W28(W28TO51), .W29(W29TO51), .W30(W30TO51), .W31(W31TO51), .W32(W32TO51), .W33(W33TO51), .W34(W34TO51), .W35(W35TO51), .W36(W36TO51), .W37(W37TO51), .W38(W38TO51), .W39(W39TO51), .W40(W40TO51), .W41(W41TO51), .W42(W42TO51), .W43(W43TO51), .W44(W44TO51), .W45(W45TO51), .W46(W46TO51), .W47(W47TO51), .W48(W48TO51), .W49(W49TO51), .W50(W50TO51), .W51(W51TO51), .W52(W52TO51), .W53(W53TO51), .W54(W54TO51), .W55(W55TO51), .W56(W56TO51), .W57(W57TO51), .W58(W58TO51), .W59(W59TO51), .W60(W60TO51), .W61(W61TO51), .W62(W62TO51), .W63(W63TO51)) neuron51(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out51));
neuron64in #(.W0(W0TO52), .W1(W1TO52), .W2(W2TO52), .W3(W3TO52), .W4(W4TO52), .W5(W5TO52), .W6(W6TO52), .W7(W7TO52), .W8(W8TO52), .W9(W9TO52), .W10(W10TO52), .W11(W11TO52), .W12(W12TO52), .W13(W13TO52), .W14(W14TO52), .W15(W15TO52), .W16(W16TO52), .W17(W17TO52), .W18(W18TO52), .W19(W19TO52), .W20(W20TO52), .W21(W21TO52), .W22(W22TO52), .W23(W23TO52), .W24(W24TO52), .W25(W25TO52), .W26(W26TO52), .W27(W27TO52), .W28(W28TO52), .W29(W29TO52), .W30(W30TO52), .W31(W31TO52), .W32(W32TO52), .W33(W33TO52), .W34(W34TO52), .W35(W35TO52), .W36(W36TO52), .W37(W37TO52), .W38(W38TO52), .W39(W39TO52), .W40(W40TO52), .W41(W41TO52), .W42(W42TO52), .W43(W43TO52), .W44(W44TO52), .W45(W45TO52), .W46(W46TO52), .W47(W47TO52), .W48(W48TO52), .W49(W49TO52), .W50(W50TO52), .W51(W51TO52), .W52(W52TO52), .W53(W53TO52), .W54(W54TO52), .W55(W55TO52), .W56(W56TO52), .W57(W57TO52), .W58(W58TO52), .W59(W59TO52), .W60(W60TO52), .W61(W61TO52), .W62(W62TO52), .W63(W63TO52)) neuron52(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out52));
neuron64in #(.W0(W0TO53), .W1(W1TO53), .W2(W2TO53), .W3(W3TO53), .W4(W4TO53), .W5(W5TO53), .W6(W6TO53), .W7(W7TO53), .W8(W8TO53), .W9(W9TO53), .W10(W10TO53), .W11(W11TO53), .W12(W12TO53), .W13(W13TO53), .W14(W14TO53), .W15(W15TO53), .W16(W16TO53), .W17(W17TO53), .W18(W18TO53), .W19(W19TO53), .W20(W20TO53), .W21(W21TO53), .W22(W22TO53), .W23(W23TO53), .W24(W24TO53), .W25(W25TO53), .W26(W26TO53), .W27(W27TO53), .W28(W28TO53), .W29(W29TO53), .W30(W30TO53), .W31(W31TO53), .W32(W32TO53), .W33(W33TO53), .W34(W34TO53), .W35(W35TO53), .W36(W36TO53), .W37(W37TO53), .W38(W38TO53), .W39(W39TO53), .W40(W40TO53), .W41(W41TO53), .W42(W42TO53), .W43(W43TO53), .W44(W44TO53), .W45(W45TO53), .W46(W46TO53), .W47(W47TO53), .W48(W48TO53), .W49(W49TO53), .W50(W50TO53), .W51(W51TO53), .W52(W52TO53), .W53(W53TO53), .W54(W54TO53), .W55(W55TO53), .W56(W56TO53), .W57(W57TO53), .W58(W58TO53), .W59(W59TO53), .W60(W60TO53), .W61(W61TO53), .W62(W62TO53), .W63(W63TO53)) neuron53(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out53));
neuron64in #(.W0(W0TO54), .W1(W1TO54), .W2(W2TO54), .W3(W3TO54), .W4(W4TO54), .W5(W5TO54), .W6(W6TO54), .W7(W7TO54), .W8(W8TO54), .W9(W9TO54), .W10(W10TO54), .W11(W11TO54), .W12(W12TO54), .W13(W13TO54), .W14(W14TO54), .W15(W15TO54), .W16(W16TO54), .W17(W17TO54), .W18(W18TO54), .W19(W19TO54), .W20(W20TO54), .W21(W21TO54), .W22(W22TO54), .W23(W23TO54), .W24(W24TO54), .W25(W25TO54), .W26(W26TO54), .W27(W27TO54), .W28(W28TO54), .W29(W29TO54), .W30(W30TO54), .W31(W31TO54), .W32(W32TO54), .W33(W33TO54), .W34(W34TO54), .W35(W35TO54), .W36(W36TO54), .W37(W37TO54), .W38(W38TO54), .W39(W39TO54), .W40(W40TO54), .W41(W41TO54), .W42(W42TO54), .W43(W43TO54), .W44(W44TO54), .W45(W45TO54), .W46(W46TO54), .W47(W47TO54), .W48(W48TO54), .W49(W49TO54), .W50(W50TO54), .W51(W51TO54), .W52(W52TO54), .W53(W53TO54), .W54(W54TO54), .W55(W55TO54), .W56(W56TO54), .W57(W57TO54), .W58(W58TO54), .W59(W59TO54), .W60(W60TO54), .W61(W61TO54), .W62(W62TO54), .W63(W63TO54)) neuron54(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out54));
neuron64in #(.W0(W0TO55), .W1(W1TO55), .W2(W2TO55), .W3(W3TO55), .W4(W4TO55), .W5(W5TO55), .W6(W6TO55), .W7(W7TO55), .W8(W8TO55), .W9(W9TO55), .W10(W10TO55), .W11(W11TO55), .W12(W12TO55), .W13(W13TO55), .W14(W14TO55), .W15(W15TO55), .W16(W16TO55), .W17(W17TO55), .W18(W18TO55), .W19(W19TO55), .W20(W20TO55), .W21(W21TO55), .W22(W22TO55), .W23(W23TO55), .W24(W24TO55), .W25(W25TO55), .W26(W26TO55), .W27(W27TO55), .W28(W28TO55), .W29(W29TO55), .W30(W30TO55), .W31(W31TO55), .W32(W32TO55), .W33(W33TO55), .W34(W34TO55), .W35(W35TO55), .W36(W36TO55), .W37(W37TO55), .W38(W38TO55), .W39(W39TO55), .W40(W40TO55), .W41(W41TO55), .W42(W42TO55), .W43(W43TO55), .W44(W44TO55), .W45(W45TO55), .W46(W46TO55), .W47(W47TO55), .W48(W48TO55), .W49(W49TO55), .W50(W50TO55), .W51(W51TO55), .W52(W52TO55), .W53(W53TO55), .W54(W54TO55), .W55(W55TO55), .W56(W56TO55), .W57(W57TO55), .W58(W58TO55), .W59(W59TO55), .W60(W60TO55), .W61(W61TO55), .W62(W62TO55), .W63(W63TO55)) neuron55(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out55));
neuron64in #(.W0(W0TO56), .W1(W1TO56), .W2(W2TO56), .W3(W3TO56), .W4(W4TO56), .W5(W5TO56), .W6(W6TO56), .W7(W7TO56), .W8(W8TO56), .W9(W9TO56), .W10(W10TO56), .W11(W11TO56), .W12(W12TO56), .W13(W13TO56), .W14(W14TO56), .W15(W15TO56), .W16(W16TO56), .W17(W17TO56), .W18(W18TO56), .W19(W19TO56), .W20(W20TO56), .W21(W21TO56), .W22(W22TO56), .W23(W23TO56), .W24(W24TO56), .W25(W25TO56), .W26(W26TO56), .W27(W27TO56), .W28(W28TO56), .W29(W29TO56), .W30(W30TO56), .W31(W31TO56), .W32(W32TO56), .W33(W33TO56), .W34(W34TO56), .W35(W35TO56), .W36(W36TO56), .W37(W37TO56), .W38(W38TO56), .W39(W39TO56), .W40(W40TO56), .W41(W41TO56), .W42(W42TO56), .W43(W43TO56), .W44(W44TO56), .W45(W45TO56), .W46(W46TO56), .W47(W47TO56), .W48(W48TO56), .W49(W49TO56), .W50(W50TO56), .W51(W51TO56), .W52(W52TO56), .W53(W53TO56), .W54(W54TO56), .W55(W55TO56), .W56(W56TO56), .W57(W57TO56), .W58(W58TO56), .W59(W59TO56), .W60(W60TO56), .W61(W61TO56), .W62(W62TO56), .W63(W63TO56)) neuron56(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out56));
neuron64in #(.W0(W0TO57), .W1(W1TO57), .W2(W2TO57), .W3(W3TO57), .W4(W4TO57), .W5(W5TO57), .W6(W6TO57), .W7(W7TO57), .W8(W8TO57), .W9(W9TO57), .W10(W10TO57), .W11(W11TO57), .W12(W12TO57), .W13(W13TO57), .W14(W14TO57), .W15(W15TO57), .W16(W16TO57), .W17(W17TO57), .W18(W18TO57), .W19(W19TO57), .W20(W20TO57), .W21(W21TO57), .W22(W22TO57), .W23(W23TO57), .W24(W24TO57), .W25(W25TO57), .W26(W26TO57), .W27(W27TO57), .W28(W28TO57), .W29(W29TO57), .W30(W30TO57), .W31(W31TO57), .W32(W32TO57), .W33(W33TO57), .W34(W34TO57), .W35(W35TO57), .W36(W36TO57), .W37(W37TO57), .W38(W38TO57), .W39(W39TO57), .W40(W40TO57), .W41(W41TO57), .W42(W42TO57), .W43(W43TO57), .W44(W44TO57), .W45(W45TO57), .W46(W46TO57), .W47(W47TO57), .W48(W48TO57), .W49(W49TO57), .W50(W50TO57), .W51(W51TO57), .W52(W52TO57), .W53(W53TO57), .W54(W54TO57), .W55(W55TO57), .W56(W56TO57), .W57(W57TO57), .W58(W58TO57), .W59(W59TO57), .W60(W60TO57), .W61(W61TO57), .W62(W62TO57), .W63(W63TO57)) neuron57(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out57));
neuron64in #(.W0(W0TO58), .W1(W1TO58), .W2(W2TO58), .W3(W3TO58), .W4(W4TO58), .W5(W5TO58), .W6(W6TO58), .W7(W7TO58), .W8(W8TO58), .W9(W9TO58), .W10(W10TO58), .W11(W11TO58), .W12(W12TO58), .W13(W13TO58), .W14(W14TO58), .W15(W15TO58), .W16(W16TO58), .W17(W17TO58), .W18(W18TO58), .W19(W19TO58), .W20(W20TO58), .W21(W21TO58), .W22(W22TO58), .W23(W23TO58), .W24(W24TO58), .W25(W25TO58), .W26(W26TO58), .W27(W27TO58), .W28(W28TO58), .W29(W29TO58), .W30(W30TO58), .W31(W31TO58), .W32(W32TO58), .W33(W33TO58), .W34(W34TO58), .W35(W35TO58), .W36(W36TO58), .W37(W37TO58), .W38(W38TO58), .W39(W39TO58), .W40(W40TO58), .W41(W41TO58), .W42(W42TO58), .W43(W43TO58), .W44(W44TO58), .W45(W45TO58), .W46(W46TO58), .W47(W47TO58), .W48(W48TO58), .W49(W49TO58), .W50(W50TO58), .W51(W51TO58), .W52(W52TO58), .W53(W53TO58), .W54(W54TO58), .W55(W55TO58), .W56(W56TO58), .W57(W57TO58), .W58(W58TO58), .W59(W59TO58), .W60(W60TO58), .W61(W61TO58), .W62(W62TO58), .W63(W63TO58)) neuron58(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out58));
neuron64in #(.W0(W0TO59), .W1(W1TO59), .W2(W2TO59), .W3(W3TO59), .W4(W4TO59), .W5(W5TO59), .W6(W6TO59), .W7(W7TO59), .W8(W8TO59), .W9(W9TO59), .W10(W10TO59), .W11(W11TO59), .W12(W12TO59), .W13(W13TO59), .W14(W14TO59), .W15(W15TO59), .W16(W16TO59), .W17(W17TO59), .W18(W18TO59), .W19(W19TO59), .W20(W20TO59), .W21(W21TO59), .W22(W22TO59), .W23(W23TO59), .W24(W24TO59), .W25(W25TO59), .W26(W26TO59), .W27(W27TO59), .W28(W28TO59), .W29(W29TO59), .W30(W30TO59), .W31(W31TO59), .W32(W32TO59), .W33(W33TO59), .W34(W34TO59), .W35(W35TO59), .W36(W36TO59), .W37(W37TO59), .W38(W38TO59), .W39(W39TO59), .W40(W40TO59), .W41(W41TO59), .W42(W42TO59), .W43(W43TO59), .W44(W44TO59), .W45(W45TO59), .W46(W46TO59), .W47(W47TO59), .W48(W48TO59), .W49(W49TO59), .W50(W50TO59), .W51(W51TO59), .W52(W52TO59), .W53(W53TO59), .W54(W54TO59), .W55(W55TO59), .W56(W56TO59), .W57(W57TO59), .W58(W58TO59), .W59(W59TO59), .W60(W60TO59), .W61(W61TO59), .W62(W62TO59), .W63(W63TO59)) neuron59(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out59));
neuron64in #(.W0(W0TO60), .W1(W1TO60), .W2(W2TO60), .W3(W3TO60), .W4(W4TO60), .W5(W5TO60), .W6(W6TO60), .W7(W7TO60), .W8(W8TO60), .W9(W9TO60), .W10(W10TO60), .W11(W11TO60), .W12(W12TO60), .W13(W13TO60), .W14(W14TO60), .W15(W15TO60), .W16(W16TO60), .W17(W17TO60), .W18(W18TO60), .W19(W19TO60), .W20(W20TO60), .W21(W21TO60), .W22(W22TO60), .W23(W23TO60), .W24(W24TO60), .W25(W25TO60), .W26(W26TO60), .W27(W27TO60), .W28(W28TO60), .W29(W29TO60), .W30(W30TO60), .W31(W31TO60), .W32(W32TO60), .W33(W33TO60), .W34(W34TO60), .W35(W35TO60), .W36(W36TO60), .W37(W37TO60), .W38(W38TO60), .W39(W39TO60), .W40(W40TO60), .W41(W41TO60), .W42(W42TO60), .W43(W43TO60), .W44(W44TO60), .W45(W45TO60), .W46(W46TO60), .W47(W47TO60), .W48(W48TO60), .W49(W49TO60), .W50(W50TO60), .W51(W51TO60), .W52(W52TO60), .W53(W53TO60), .W54(W54TO60), .W55(W55TO60), .W56(W56TO60), .W57(W57TO60), .W58(W58TO60), .W59(W59TO60), .W60(W60TO60), .W61(W61TO60), .W62(W62TO60), .W63(W63TO60)) neuron60(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out60));
neuron64in #(.W0(W0TO61), .W1(W1TO61), .W2(W2TO61), .W3(W3TO61), .W4(W4TO61), .W5(W5TO61), .W6(W6TO61), .W7(W7TO61), .W8(W8TO61), .W9(W9TO61), .W10(W10TO61), .W11(W11TO61), .W12(W12TO61), .W13(W13TO61), .W14(W14TO61), .W15(W15TO61), .W16(W16TO61), .W17(W17TO61), .W18(W18TO61), .W19(W19TO61), .W20(W20TO61), .W21(W21TO61), .W22(W22TO61), .W23(W23TO61), .W24(W24TO61), .W25(W25TO61), .W26(W26TO61), .W27(W27TO61), .W28(W28TO61), .W29(W29TO61), .W30(W30TO61), .W31(W31TO61), .W32(W32TO61), .W33(W33TO61), .W34(W34TO61), .W35(W35TO61), .W36(W36TO61), .W37(W37TO61), .W38(W38TO61), .W39(W39TO61), .W40(W40TO61), .W41(W41TO61), .W42(W42TO61), .W43(W43TO61), .W44(W44TO61), .W45(W45TO61), .W46(W46TO61), .W47(W47TO61), .W48(W48TO61), .W49(W49TO61), .W50(W50TO61), .W51(W51TO61), .W52(W52TO61), .W53(W53TO61), .W54(W54TO61), .W55(W55TO61), .W56(W56TO61), .W57(W57TO61), .W58(W58TO61), .W59(W59TO61), .W60(W60TO61), .W61(W61TO61), .W62(W62TO61), .W63(W63TO61)) neuron61(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out61));
neuron64in #(.W0(W0TO62), .W1(W1TO62), .W2(W2TO62), .W3(W3TO62), .W4(W4TO62), .W5(W5TO62), .W6(W6TO62), .W7(W7TO62), .W8(W8TO62), .W9(W9TO62), .W10(W10TO62), .W11(W11TO62), .W12(W12TO62), .W13(W13TO62), .W14(W14TO62), .W15(W15TO62), .W16(W16TO62), .W17(W17TO62), .W18(W18TO62), .W19(W19TO62), .W20(W20TO62), .W21(W21TO62), .W22(W22TO62), .W23(W23TO62), .W24(W24TO62), .W25(W25TO62), .W26(W26TO62), .W27(W27TO62), .W28(W28TO62), .W29(W29TO62), .W30(W30TO62), .W31(W31TO62), .W32(W32TO62), .W33(W33TO62), .W34(W34TO62), .W35(W35TO62), .W36(W36TO62), .W37(W37TO62), .W38(W38TO62), .W39(W39TO62), .W40(W40TO62), .W41(W41TO62), .W42(W42TO62), .W43(W43TO62), .W44(W44TO62), .W45(W45TO62), .W46(W46TO62), .W47(W47TO62), .W48(W48TO62), .W49(W49TO62), .W50(W50TO62), .W51(W51TO62), .W52(W52TO62), .W53(W53TO62), .W54(W54TO62), .W55(W55TO62), .W56(W56TO62), .W57(W57TO62), .W58(W58TO62), .W59(W59TO62), .W60(W60TO62), .W61(W61TO62), .W62(W62TO62), .W63(W63TO62)) neuron62(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out62));
neuron64in #(.W0(W0TO63), .W1(W1TO63), .W2(W2TO63), .W3(W3TO63), .W4(W4TO63), .W5(W5TO63), .W6(W6TO63), .W7(W7TO63), .W8(W8TO63), .W9(W9TO63), .W10(W10TO63), .W11(W11TO63), .W12(W12TO63), .W13(W13TO63), .W14(W14TO63), .W15(W15TO63), .W16(W16TO63), .W17(W17TO63), .W18(W18TO63), .W19(W19TO63), .W20(W20TO63), .W21(W21TO63), .W22(W22TO63), .W23(W23TO63), .W24(W24TO63), .W25(W25TO63), .W26(W26TO63), .W27(W27TO63), .W28(W28TO63), .W29(W29TO63), .W30(W30TO63), .W31(W31TO63), .W32(W32TO63), .W33(W33TO63), .W34(W34TO63), .W35(W35TO63), .W36(W36TO63), .W37(W37TO63), .W38(W38TO63), .W39(W39TO63), .W40(W40TO63), .W41(W41TO63), .W42(W42TO63), .W43(W43TO63), .W44(W44TO63), .W45(W45TO63), .W46(W46TO63), .W47(W47TO63), .W48(W48TO63), .W49(W49TO63), .W50(W50TO63), .W51(W51TO63), .W52(W52TO63), .W53(W53TO63), .W54(W54TO63), .W55(W55TO63), .W56(W56TO63), .W57(W57TO63), .W58(W58TO63), .W59(W59TO63), .W60(W60TO63), .W61(W61TO63), .W62(W62TO63), .W63(W63TO63)) neuron63(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out63));
neuron64in #(.W0(W0TO64), .W1(W1TO64), .W2(W2TO64), .W3(W3TO64), .W4(W4TO64), .W5(W5TO64), .W6(W6TO64), .W7(W7TO64), .W8(W8TO64), .W9(W9TO64), .W10(W10TO64), .W11(W11TO64), .W12(W12TO64), .W13(W13TO64), .W14(W14TO64), .W15(W15TO64), .W16(W16TO64), .W17(W17TO64), .W18(W18TO64), .W19(W19TO64), .W20(W20TO64), .W21(W21TO64), .W22(W22TO64), .W23(W23TO64), .W24(W24TO64), .W25(W25TO64), .W26(W26TO64), .W27(W27TO64), .W28(W28TO64), .W29(W29TO64), .W30(W30TO64), .W31(W31TO64), .W32(W32TO64), .W33(W33TO64), .W34(W34TO64), .W35(W35TO64), .W36(W36TO64), .W37(W37TO64), .W38(W38TO64), .W39(W39TO64), .W40(W40TO64), .W41(W41TO64), .W42(W42TO64), .W43(W43TO64), .W44(W44TO64), .W45(W45TO64), .W46(W46TO64), .W47(W47TO64), .W48(W48TO64), .W49(W49TO64), .W50(W50TO64), .W51(W51TO64), .W52(W52TO64), .W53(W53TO64), .W54(W54TO64), .W55(W55TO64), .W56(W56TO64), .W57(W57TO64), .W58(W58TO64), .W59(W59TO64), .W60(W60TO64), .W61(W61TO64), .W62(W62TO64), .W63(W63TO64)) neuron64(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out64));
neuron64in #(.W0(W0TO65), .W1(W1TO65), .W2(W2TO65), .W3(W3TO65), .W4(W4TO65), .W5(W5TO65), .W6(W6TO65), .W7(W7TO65), .W8(W8TO65), .W9(W9TO65), .W10(W10TO65), .W11(W11TO65), .W12(W12TO65), .W13(W13TO65), .W14(W14TO65), .W15(W15TO65), .W16(W16TO65), .W17(W17TO65), .W18(W18TO65), .W19(W19TO65), .W20(W20TO65), .W21(W21TO65), .W22(W22TO65), .W23(W23TO65), .W24(W24TO65), .W25(W25TO65), .W26(W26TO65), .W27(W27TO65), .W28(W28TO65), .W29(W29TO65), .W30(W30TO65), .W31(W31TO65), .W32(W32TO65), .W33(W33TO65), .W34(W34TO65), .W35(W35TO65), .W36(W36TO65), .W37(W37TO65), .W38(W38TO65), .W39(W39TO65), .W40(W40TO65), .W41(W41TO65), .W42(W42TO65), .W43(W43TO65), .W44(W44TO65), .W45(W45TO65), .W46(W46TO65), .W47(W47TO65), .W48(W48TO65), .W49(W49TO65), .W50(W50TO65), .W51(W51TO65), .W52(W52TO65), .W53(W53TO65), .W54(W54TO65), .W55(W55TO65), .W56(W56TO65), .W57(W57TO65), .W58(W58TO65), .W59(W59TO65), .W60(W60TO65), .W61(W61TO65), .W62(W62TO65), .W63(W63TO65)) neuron65(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out65));
neuron64in #(.W0(W0TO66), .W1(W1TO66), .W2(W2TO66), .W3(W3TO66), .W4(W4TO66), .W5(W5TO66), .W6(W6TO66), .W7(W7TO66), .W8(W8TO66), .W9(W9TO66), .W10(W10TO66), .W11(W11TO66), .W12(W12TO66), .W13(W13TO66), .W14(W14TO66), .W15(W15TO66), .W16(W16TO66), .W17(W17TO66), .W18(W18TO66), .W19(W19TO66), .W20(W20TO66), .W21(W21TO66), .W22(W22TO66), .W23(W23TO66), .W24(W24TO66), .W25(W25TO66), .W26(W26TO66), .W27(W27TO66), .W28(W28TO66), .W29(W29TO66), .W30(W30TO66), .W31(W31TO66), .W32(W32TO66), .W33(W33TO66), .W34(W34TO66), .W35(W35TO66), .W36(W36TO66), .W37(W37TO66), .W38(W38TO66), .W39(W39TO66), .W40(W40TO66), .W41(W41TO66), .W42(W42TO66), .W43(W43TO66), .W44(W44TO66), .W45(W45TO66), .W46(W46TO66), .W47(W47TO66), .W48(W48TO66), .W49(W49TO66), .W50(W50TO66), .W51(W51TO66), .W52(W52TO66), .W53(W53TO66), .W54(W54TO66), .W55(W55TO66), .W56(W56TO66), .W57(W57TO66), .W58(W58TO66), .W59(W59TO66), .W60(W60TO66), .W61(W61TO66), .W62(W62TO66), .W63(W63TO66)) neuron66(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out66));
neuron64in #(.W0(W0TO67), .W1(W1TO67), .W2(W2TO67), .W3(W3TO67), .W4(W4TO67), .W5(W5TO67), .W6(W6TO67), .W7(W7TO67), .W8(W8TO67), .W9(W9TO67), .W10(W10TO67), .W11(W11TO67), .W12(W12TO67), .W13(W13TO67), .W14(W14TO67), .W15(W15TO67), .W16(W16TO67), .W17(W17TO67), .W18(W18TO67), .W19(W19TO67), .W20(W20TO67), .W21(W21TO67), .W22(W22TO67), .W23(W23TO67), .W24(W24TO67), .W25(W25TO67), .W26(W26TO67), .W27(W27TO67), .W28(W28TO67), .W29(W29TO67), .W30(W30TO67), .W31(W31TO67), .W32(W32TO67), .W33(W33TO67), .W34(W34TO67), .W35(W35TO67), .W36(W36TO67), .W37(W37TO67), .W38(W38TO67), .W39(W39TO67), .W40(W40TO67), .W41(W41TO67), .W42(W42TO67), .W43(W43TO67), .W44(W44TO67), .W45(W45TO67), .W46(W46TO67), .W47(W47TO67), .W48(W48TO67), .W49(W49TO67), .W50(W50TO67), .W51(W51TO67), .W52(W52TO67), .W53(W53TO67), .W54(W54TO67), .W55(W55TO67), .W56(W56TO67), .W57(W57TO67), .W58(W58TO67), .W59(W59TO67), .W60(W60TO67), .W61(W61TO67), .W62(W62TO67), .W63(W63TO67)) neuron67(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out67));
neuron64in #(.W0(W0TO68), .W1(W1TO68), .W2(W2TO68), .W3(W3TO68), .W4(W4TO68), .W5(W5TO68), .W6(W6TO68), .W7(W7TO68), .W8(W8TO68), .W9(W9TO68), .W10(W10TO68), .W11(W11TO68), .W12(W12TO68), .W13(W13TO68), .W14(W14TO68), .W15(W15TO68), .W16(W16TO68), .W17(W17TO68), .W18(W18TO68), .W19(W19TO68), .W20(W20TO68), .W21(W21TO68), .W22(W22TO68), .W23(W23TO68), .W24(W24TO68), .W25(W25TO68), .W26(W26TO68), .W27(W27TO68), .W28(W28TO68), .W29(W29TO68), .W30(W30TO68), .W31(W31TO68), .W32(W32TO68), .W33(W33TO68), .W34(W34TO68), .W35(W35TO68), .W36(W36TO68), .W37(W37TO68), .W38(W38TO68), .W39(W39TO68), .W40(W40TO68), .W41(W41TO68), .W42(W42TO68), .W43(W43TO68), .W44(W44TO68), .W45(W45TO68), .W46(W46TO68), .W47(W47TO68), .W48(W48TO68), .W49(W49TO68), .W50(W50TO68), .W51(W51TO68), .W52(W52TO68), .W53(W53TO68), .W54(W54TO68), .W55(W55TO68), .W56(W56TO68), .W57(W57TO68), .W58(W58TO68), .W59(W59TO68), .W60(W60TO68), .W61(W61TO68), .W62(W62TO68), .W63(W63TO68)) neuron68(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out68));
neuron64in #(.W0(W0TO69), .W1(W1TO69), .W2(W2TO69), .W3(W3TO69), .W4(W4TO69), .W5(W5TO69), .W6(W6TO69), .W7(W7TO69), .W8(W8TO69), .W9(W9TO69), .W10(W10TO69), .W11(W11TO69), .W12(W12TO69), .W13(W13TO69), .W14(W14TO69), .W15(W15TO69), .W16(W16TO69), .W17(W17TO69), .W18(W18TO69), .W19(W19TO69), .W20(W20TO69), .W21(W21TO69), .W22(W22TO69), .W23(W23TO69), .W24(W24TO69), .W25(W25TO69), .W26(W26TO69), .W27(W27TO69), .W28(W28TO69), .W29(W29TO69), .W30(W30TO69), .W31(W31TO69), .W32(W32TO69), .W33(W33TO69), .W34(W34TO69), .W35(W35TO69), .W36(W36TO69), .W37(W37TO69), .W38(W38TO69), .W39(W39TO69), .W40(W40TO69), .W41(W41TO69), .W42(W42TO69), .W43(W43TO69), .W44(W44TO69), .W45(W45TO69), .W46(W46TO69), .W47(W47TO69), .W48(W48TO69), .W49(W49TO69), .W50(W50TO69), .W51(W51TO69), .W52(W52TO69), .W53(W53TO69), .W54(W54TO69), .W55(W55TO69), .W56(W56TO69), .W57(W57TO69), .W58(W58TO69), .W59(W59TO69), .W60(W60TO69), .W61(W61TO69), .W62(W62TO69), .W63(W63TO69)) neuron69(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out69));
neuron64in #(.W0(W0TO70), .W1(W1TO70), .W2(W2TO70), .W3(W3TO70), .W4(W4TO70), .W5(W5TO70), .W6(W6TO70), .W7(W7TO70), .W8(W8TO70), .W9(W9TO70), .W10(W10TO70), .W11(W11TO70), .W12(W12TO70), .W13(W13TO70), .W14(W14TO70), .W15(W15TO70), .W16(W16TO70), .W17(W17TO70), .W18(W18TO70), .W19(W19TO70), .W20(W20TO70), .W21(W21TO70), .W22(W22TO70), .W23(W23TO70), .W24(W24TO70), .W25(W25TO70), .W26(W26TO70), .W27(W27TO70), .W28(W28TO70), .W29(W29TO70), .W30(W30TO70), .W31(W31TO70), .W32(W32TO70), .W33(W33TO70), .W34(W34TO70), .W35(W35TO70), .W36(W36TO70), .W37(W37TO70), .W38(W38TO70), .W39(W39TO70), .W40(W40TO70), .W41(W41TO70), .W42(W42TO70), .W43(W43TO70), .W44(W44TO70), .W45(W45TO70), .W46(W46TO70), .W47(W47TO70), .W48(W48TO70), .W49(W49TO70), .W50(W50TO70), .W51(W51TO70), .W52(W52TO70), .W53(W53TO70), .W54(W54TO70), .W55(W55TO70), .W56(W56TO70), .W57(W57TO70), .W58(W58TO70), .W59(W59TO70), .W60(W60TO70), .W61(W61TO70), .W62(W62TO70), .W63(W63TO70)) neuron70(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out70));
neuron64in #(.W0(W0TO71), .W1(W1TO71), .W2(W2TO71), .W3(W3TO71), .W4(W4TO71), .W5(W5TO71), .W6(W6TO71), .W7(W7TO71), .W8(W8TO71), .W9(W9TO71), .W10(W10TO71), .W11(W11TO71), .W12(W12TO71), .W13(W13TO71), .W14(W14TO71), .W15(W15TO71), .W16(W16TO71), .W17(W17TO71), .W18(W18TO71), .W19(W19TO71), .W20(W20TO71), .W21(W21TO71), .W22(W22TO71), .W23(W23TO71), .W24(W24TO71), .W25(W25TO71), .W26(W26TO71), .W27(W27TO71), .W28(W28TO71), .W29(W29TO71), .W30(W30TO71), .W31(W31TO71), .W32(W32TO71), .W33(W33TO71), .W34(W34TO71), .W35(W35TO71), .W36(W36TO71), .W37(W37TO71), .W38(W38TO71), .W39(W39TO71), .W40(W40TO71), .W41(W41TO71), .W42(W42TO71), .W43(W43TO71), .W44(W44TO71), .W45(W45TO71), .W46(W46TO71), .W47(W47TO71), .W48(W48TO71), .W49(W49TO71), .W50(W50TO71), .W51(W51TO71), .W52(W52TO71), .W53(W53TO71), .W54(W54TO71), .W55(W55TO71), .W56(W56TO71), .W57(W57TO71), .W58(W58TO71), .W59(W59TO71), .W60(W60TO71), .W61(W61TO71), .W62(W62TO71), .W63(W63TO71)) neuron71(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out71));
neuron64in #(.W0(W0TO72), .W1(W1TO72), .W2(W2TO72), .W3(W3TO72), .W4(W4TO72), .W5(W5TO72), .W6(W6TO72), .W7(W7TO72), .W8(W8TO72), .W9(W9TO72), .W10(W10TO72), .W11(W11TO72), .W12(W12TO72), .W13(W13TO72), .W14(W14TO72), .W15(W15TO72), .W16(W16TO72), .W17(W17TO72), .W18(W18TO72), .W19(W19TO72), .W20(W20TO72), .W21(W21TO72), .W22(W22TO72), .W23(W23TO72), .W24(W24TO72), .W25(W25TO72), .W26(W26TO72), .W27(W27TO72), .W28(W28TO72), .W29(W29TO72), .W30(W30TO72), .W31(W31TO72), .W32(W32TO72), .W33(W33TO72), .W34(W34TO72), .W35(W35TO72), .W36(W36TO72), .W37(W37TO72), .W38(W38TO72), .W39(W39TO72), .W40(W40TO72), .W41(W41TO72), .W42(W42TO72), .W43(W43TO72), .W44(W44TO72), .W45(W45TO72), .W46(W46TO72), .W47(W47TO72), .W48(W48TO72), .W49(W49TO72), .W50(W50TO72), .W51(W51TO72), .W52(W52TO72), .W53(W53TO72), .W54(W54TO72), .W55(W55TO72), .W56(W56TO72), .W57(W57TO72), .W58(W58TO72), .W59(W59TO72), .W60(W60TO72), .W61(W61TO72), .W62(W62TO72), .W63(W63TO72)) neuron72(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out72));
neuron64in #(.W0(W0TO73), .W1(W1TO73), .W2(W2TO73), .W3(W3TO73), .W4(W4TO73), .W5(W5TO73), .W6(W6TO73), .W7(W7TO73), .W8(W8TO73), .W9(W9TO73), .W10(W10TO73), .W11(W11TO73), .W12(W12TO73), .W13(W13TO73), .W14(W14TO73), .W15(W15TO73), .W16(W16TO73), .W17(W17TO73), .W18(W18TO73), .W19(W19TO73), .W20(W20TO73), .W21(W21TO73), .W22(W22TO73), .W23(W23TO73), .W24(W24TO73), .W25(W25TO73), .W26(W26TO73), .W27(W27TO73), .W28(W28TO73), .W29(W29TO73), .W30(W30TO73), .W31(W31TO73), .W32(W32TO73), .W33(W33TO73), .W34(W34TO73), .W35(W35TO73), .W36(W36TO73), .W37(W37TO73), .W38(W38TO73), .W39(W39TO73), .W40(W40TO73), .W41(W41TO73), .W42(W42TO73), .W43(W43TO73), .W44(W44TO73), .W45(W45TO73), .W46(W46TO73), .W47(W47TO73), .W48(W48TO73), .W49(W49TO73), .W50(W50TO73), .W51(W51TO73), .W52(W52TO73), .W53(W53TO73), .W54(W54TO73), .W55(W55TO73), .W56(W56TO73), .W57(W57TO73), .W58(W58TO73), .W59(W59TO73), .W60(W60TO73), .W61(W61TO73), .W62(W62TO73), .W63(W63TO73)) neuron73(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out73));
neuron64in #(.W0(W0TO74), .W1(W1TO74), .W2(W2TO74), .W3(W3TO74), .W4(W4TO74), .W5(W5TO74), .W6(W6TO74), .W7(W7TO74), .W8(W8TO74), .W9(W9TO74), .W10(W10TO74), .W11(W11TO74), .W12(W12TO74), .W13(W13TO74), .W14(W14TO74), .W15(W15TO74), .W16(W16TO74), .W17(W17TO74), .W18(W18TO74), .W19(W19TO74), .W20(W20TO74), .W21(W21TO74), .W22(W22TO74), .W23(W23TO74), .W24(W24TO74), .W25(W25TO74), .W26(W26TO74), .W27(W27TO74), .W28(W28TO74), .W29(W29TO74), .W30(W30TO74), .W31(W31TO74), .W32(W32TO74), .W33(W33TO74), .W34(W34TO74), .W35(W35TO74), .W36(W36TO74), .W37(W37TO74), .W38(W38TO74), .W39(W39TO74), .W40(W40TO74), .W41(W41TO74), .W42(W42TO74), .W43(W43TO74), .W44(W44TO74), .W45(W45TO74), .W46(W46TO74), .W47(W47TO74), .W48(W48TO74), .W49(W49TO74), .W50(W50TO74), .W51(W51TO74), .W52(W52TO74), .W53(W53TO74), .W54(W54TO74), .W55(W55TO74), .W56(W56TO74), .W57(W57TO74), .W58(W58TO74), .W59(W59TO74), .W60(W60TO74), .W61(W61TO74), .W62(W62TO74), .W63(W63TO74)) neuron74(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out74));
neuron64in #(.W0(W0TO75), .W1(W1TO75), .W2(W2TO75), .W3(W3TO75), .W4(W4TO75), .W5(W5TO75), .W6(W6TO75), .W7(W7TO75), .W8(W8TO75), .W9(W9TO75), .W10(W10TO75), .W11(W11TO75), .W12(W12TO75), .W13(W13TO75), .W14(W14TO75), .W15(W15TO75), .W16(W16TO75), .W17(W17TO75), .W18(W18TO75), .W19(W19TO75), .W20(W20TO75), .W21(W21TO75), .W22(W22TO75), .W23(W23TO75), .W24(W24TO75), .W25(W25TO75), .W26(W26TO75), .W27(W27TO75), .W28(W28TO75), .W29(W29TO75), .W30(W30TO75), .W31(W31TO75), .W32(W32TO75), .W33(W33TO75), .W34(W34TO75), .W35(W35TO75), .W36(W36TO75), .W37(W37TO75), .W38(W38TO75), .W39(W39TO75), .W40(W40TO75), .W41(W41TO75), .W42(W42TO75), .W43(W43TO75), .W44(W44TO75), .W45(W45TO75), .W46(W46TO75), .W47(W47TO75), .W48(W48TO75), .W49(W49TO75), .W50(W50TO75), .W51(W51TO75), .W52(W52TO75), .W53(W53TO75), .W54(W54TO75), .W55(W55TO75), .W56(W56TO75), .W57(W57TO75), .W58(W58TO75), .W59(W59TO75), .W60(W60TO75), .W61(W61TO75), .W62(W62TO75), .W63(W63TO75)) neuron75(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out75));
neuron64in #(.W0(W0TO76), .W1(W1TO76), .W2(W2TO76), .W3(W3TO76), .W4(W4TO76), .W5(W5TO76), .W6(W6TO76), .W7(W7TO76), .W8(W8TO76), .W9(W9TO76), .W10(W10TO76), .W11(W11TO76), .W12(W12TO76), .W13(W13TO76), .W14(W14TO76), .W15(W15TO76), .W16(W16TO76), .W17(W17TO76), .W18(W18TO76), .W19(W19TO76), .W20(W20TO76), .W21(W21TO76), .W22(W22TO76), .W23(W23TO76), .W24(W24TO76), .W25(W25TO76), .W26(W26TO76), .W27(W27TO76), .W28(W28TO76), .W29(W29TO76), .W30(W30TO76), .W31(W31TO76), .W32(W32TO76), .W33(W33TO76), .W34(W34TO76), .W35(W35TO76), .W36(W36TO76), .W37(W37TO76), .W38(W38TO76), .W39(W39TO76), .W40(W40TO76), .W41(W41TO76), .W42(W42TO76), .W43(W43TO76), .W44(W44TO76), .W45(W45TO76), .W46(W46TO76), .W47(W47TO76), .W48(W48TO76), .W49(W49TO76), .W50(W50TO76), .W51(W51TO76), .W52(W52TO76), .W53(W53TO76), .W54(W54TO76), .W55(W55TO76), .W56(W56TO76), .W57(W57TO76), .W58(W58TO76), .W59(W59TO76), .W60(W60TO76), .W61(W61TO76), .W62(W62TO76), .W63(W63TO76)) neuron76(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out76));
neuron64in #(.W0(W0TO77), .W1(W1TO77), .W2(W2TO77), .W3(W3TO77), .W4(W4TO77), .W5(W5TO77), .W6(W6TO77), .W7(W7TO77), .W8(W8TO77), .W9(W9TO77), .W10(W10TO77), .W11(W11TO77), .W12(W12TO77), .W13(W13TO77), .W14(W14TO77), .W15(W15TO77), .W16(W16TO77), .W17(W17TO77), .W18(W18TO77), .W19(W19TO77), .W20(W20TO77), .W21(W21TO77), .W22(W22TO77), .W23(W23TO77), .W24(W24TO77), .W25(W25TO77), .W26(W26TO77), .W27(W27TO77), .W28(W28TO77), .W29(W29TO77), .W30(W30TO77), .W31(W31TO77), .W32(W32TO77), .W33(W33TO77), .W34(W34TO77), .W35(W35TO77), .W36(W36TO77), .W37(W37TO77), .W38(W38TO77), .W39(W39TO77), .W40(W40TO77), .W41(W41TO77), .W42(W42TO77), .W43(W43TO77), .W44(W44TO77), .W45(W45TO77), .W46(W46TO77), .W47(W47TO77), .W48(W48TO77), .W49(W49TO77), .W50(W50TO77), .W51(W51TO77), .W52(W52TO77), .W53(W53TO77), .W54(W54TO77), .W55(W55TO77), .W56(W56TO77), .W57(W57TO77), .W58(W58TO77), .W59(W59TO77), .W60(W60TO77), .W61(W61TO77), .W62(W62TO77), .W63(W63TO77)) neuron77(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out77));
neuron64in #(.W0(W0TO78), .W1(W1TO78), .W2(W2TO78), .W3(W3TO78), .W4(W4TO78), .W5(W5TO78), .W6(W6TO78), .W7(W7TO78), .W8(W8TO78), .W9(W9TO78), .W10(W10TO78), .W11(W11TO78), .W12(W12TO78), .W13(W13TO78), .W14(W14TO78), .W15(W15TO78), .W16(W16TO78), .W17(W17TO78), .W18(W18TO78), .W19(W19TO78), .W20(W20TO78), .W21(W21TO78), .W22(W22TO78), .W23(W23TO78), .W24(W24TO78), .W25(W25TO78), .W26(W26TO78), .W27(W27TO78), .W28(W28TO78), .W29(W29TO78), .W30(W30TO78), .W31(W31TO78), .W32(W32TO78), .W33(W33TO78), .W34(W34TO78), .W35(W35TO78), .W36(W36TO78), .W37(W37TO78), .W38(W38TO78), .W39(W39TO78), .W40(W40TO78), .W41(W41TO78), .W42(W42TO78), .W43(W43TO78), .W44(W44TO78), .W45(W45TO78), .W46(W46TO78), .W47(W47TO78), .W48(W48TO78), .W49(W49TO78), .W50(W50TO78), .W51(W51TO78), .W52(W52TO78), .W53(W53TO78), .W54(W54TO78), .W55(W55TO78), .W56(W56TO78), .W57(W57TO78), .W58(W58TO78), .W59(W59TO78), .W60(W60TO78), .W61(W61TO78), .W62(W62TO78), .W63(W63TO78)) neuron78(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out78));
neuron64in #(.W0(W0TO79), .W1(W1TO79), .W2(W2TO79), .W3(W3TO79), .W4(W4TO79), .W5(W5TO79), .W6(W6TO79), .W7(W7TO79), .W8(W8TO79), .W9(W9TO79), .W10(W10TO79), .W11(W11TO79), .W12(W12TO79), .W13(W13TO79), .W14(W14TO79), .W15(W15TO79), .W16(W16TO79), .W17(W17TO79), .W18(W18TO79), .W19(W19TO79), .W20(W20TO79), .W21(W21TO79), .W22(W22TO79), .W23(W23TO79), .W24(W24TO79), .W25(W25TO79), .W26(W26TO79), .W27(W27TO79), .W28(W28TO79), .W29(W29TO79), .W30(W30TO79), .W31(W31TO79), .W32(W32TO79), .W33(W33TO79), .W34(W34TO79), .W35(W35TO79), .W36(W36TO79), .W37(W37TO79), .W38(W38TO79), .W39(W39TO79), .W40(W40TO79), .W41(W41TO79), .W42(W42TO79), .W43(W43TO79), .W44(W44TO79), .W45(W45TO79), .W46(W46TO79), .W47(W47TO79), .W48(W48TO79), .W49(W49TO79), .W50(W50TO79), .W51(W51TO79), .W52(W52TO79), .W53(W53TO79), .W54(W54TO79), .W55(W55TO79), .W56(W56TO79), .W57(W57TO79), .W58(W58TO79), .W59(W59TO79), .W60(W60TO79), .W61(W61TO79), .W62(W62TO79), .W63(W63TO79)) neuron79(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out79));
neuron64in #(.W0(W0TO80), .W1(W1TO80), .W2(W2TO80), .W3(W3TO80), .W4(W4TO80), .W5(W5TO80), .W6(W6TO80), .W7(W7TO80), .W8(W8TO80), .W9(W9TO80), .W10(W10TO80), .W11(W11TO80), .W12(W12TO80), .W13(W13TO80), .W14(W14TO80), .W15(W15TO80), .W16(W16TO80), .W17(W17TO80), .W18(W18TO80), .W19(W19TO80), .W20(W20TO80), .W21(W21TO80), .W22(W22TO80), .W23(W23TO80), .W24(W24TO80), .W25(W25TO80), .W26(W26TO80), .W27(W27TO80), .W28(W28TO80), .W29(W29TO80), .W30(W30TO80), .W31(W31TO80), .W32(W32TO80), .W33(W33TO80), .W34(W34TO80), .W35(W35TO80), .W36(W36TO80), .W37(W37TO80), .W38(W38TO80), .W39(W39TO80), .W40(W40TO80), .W41(W41TO80), .W42(W42TO80), .W43(W43TO80), .W44(W44TO80), .W45(W45TO80), .W46(W46TO80), .W47(W47TO80), .W48(W48TO80), .W49(W49TO80), .W50(W50TO80), .W51(W51TO80), .W52(W52TO80), .W53(W53TO80), .W54(W54TO80), .W55(W55TO80), .W56(W56TO80), .W57(W57TO80), .W58(W58TO80), .W59(W59TO80), .W60(W60TO80), .W61(W61TO80), .W62(W62TO80), .W63(W63TO80)) neuron80(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out80));
neuron64in #(.W0(W0TO81), .W1(W1TO81), .W2(W2TO81), .W3(W3TO81), .W4(W4TO81), .W5(W5TO81), .W6(W6TO81), .W7(W7TO81), .W8(W8TO81), .W9(W9TO81), .W10(W10TO81), .W11(W11TO81), .W12(W12TO81), .W13(W13TO81), .W14(W14TO81), .W15(W15TO81), .W16(W16TO81), .W17(W17TO81), .W18(W18TO81), .W19(W19TO81), .W20(W20TO81), .W21(W21TO81), .W22(W22TO81), .W23(W23TO81), .W24(W24TO81), .W25(W25TO81), .W26(W26TO81), .W27(W27TO81), .W28(W28TO81), .W29(W29TO81), .W30(W30TO81), .W31(W31TO81), .W32(W32TO81), .W33(W33TO81), .W34(W34TO81), .W35(W35TO81), .W36(W36TO81), .W37(W37TO81), .W38(W38TO81), .W39(W39TO81), .W40(W40TO81), .W41(W41TO81), .W42(W42TO81), .W43(W43TO81), .W44(W44TO81), .W45(W45TO81), .W46(W46TO81), .W47(W47TO81), .W48(W48TO81), .W49(W49TO81), .W50(W50TO81), .W51(W51TO81), .W52(W52TO81), .W53(W53TO81), .W54(W54TO81), .W55(W55TO81), .W56(W56TO81), .W57(W57TO81), .W58(W58TO81), .W59(W59TO81), .W60(W60TO81), .W61(W61TO81), .W62(W62TO81), .W63(W63TO81)) neuron81(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out81));
neuron64in #(.W0(W0TO82), .W1(W1TO82), .W2(W2TO82), .W3(W3TO82), .W4(W4TO82), .W5(W5TO82), .W6(W6TO82), .W7(W7TO82), .W8(W8TO82), .W9(W9TO82), .W10(W10TO82), .W11(W11TO82), .W12(W12TO82), .W13(W13TO82), .W14(W14TO82), .W15(W15TO82), .W16(W16TO82), .W17(W17TO82), .W18(W18TO82), .W19(W19TO82), .W20(W20TO82), .W21(W21TO82), .W22(W22TO82), .W23(W23TO82), .W24(W24TO82), .W25(W25TO82), .W26(W26TO82), .W27(W27TO82), .W28(W28TO82), .W29(W29TO82), .W30(W30TO82), .W31(W31TO82), .W32(W32TO82), .W33(W33TO82), .W34(W34TO82), .W35(W35TO82), .W36(W36TO82), .W37(W37TO82), .W38(W38TO82), .W39(W39TO82), .W40(W40TO82), .W41(W41TO82), .W42(W42TO82), .W43(W43TO82), .W44(W44TO82), .W45(W45TO82), .W46(W46TO82), .W47(W47TO82), .W48(W48TO82), .W49(W49TO82), .W50(W50TO82), .W51(W51TO82), .W52(W52TO82), .W53(W53TO82), .W54(W54TO82), .W55(W55TO82), .W56(W56TO82), .W57(W57TO82), .W58(W58TO82), .W59(W59TO82), .W60(W60TO82), .W61(W61TO82), .W62(W62TO82), .W63(W63TO82)) neuron82(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out82));
neuron64in #(.W0(W0TO83), .W1(W1TO83), .W2(W2TO83), .W3(W3TO83), .W4(W4TO83), .W5(W5TO83), .W6(W6TO83), .W7(W7TO83), .W8(W8TO83), .W9(W9TO83), .W10(W10TO83), .W11(W11TO83), .W12(W12TO83), .W13(W13TO83), .W14(W14TO83), .W15(W15TO83), .W16(W16TO83), .W17(W17TO83), .W18(W18TO83), .W19(W19TO83), .W20(W20TO83), .W21(W21TO83), .W22(W22TO83), .W23(W23TO83), .W24(W24TO83), .W25(W25TO83), .W26(W26TO83), .W27(W27TO83), .W28(W28TO83), .W29(W29TO83), .W30(W30TO83), .W31(W31TO83), .W32(W32TO83), .W33(W33TO83), .W34(W34TO83), .W35(W35TO83), .W36(W36TO83), .W37(W37TO83), .W38(W38TO83), .W39(W39TO83), .W40(W40TO83), .W41(W41TO83), .W42(W42TO83), .W43(W43TO83), .W44(W44TO83), .W45(W45TO83), .W46(W46TO83), .W47(W47TO83), .W48(W48TO83), .W49(W49TO83), .W50(W50TO83), .W51(W51TO83), .W52(W52TO83), .W53(W53TO83), .W54(W54TO83), .W55(W55TO83), .W56(W56TO83), .W57(W57TO83), .W58(W58TO83), .W59(W59TO83), .W60(W60TO83), .W61(W61TO83), .W62(W62TO83), .W63(W63TO83)) neuron83(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out83));
neuron64in #(.W0(W0TO84), .W1(W1TO84), .W2(W2TO84), .W3(W3TO84), .W4(W4TO84), .W5(W5TO84), .W6(W6TO84), .W7(W7TO84), .W8(W8TO84), .W9(W9TO84), .W10(W10TO84), .W11(W11TO84), .W12(W12TO84), .W13(W13TO84), .W14(W14TO84), .W15(W15TO84), .W16(W16TO84), .W17(W17TO84), .W18(W18TO84), .W19(W19TO84), .W20(W20TO84), .W21(W21TO84), .W22(W22TO84), .W23(W23TO84), .W24(W24TO84), .W25(W25TO84), .W26(W26TO84), .W27(W27TO84), .W28(W28TO84), .W29(W29TO84), .W30(W30TO84), .W31(W31TO84), .W32(W32TO84), .W33(W33TO84), .W34(W34TO84), .W35(W35TO84), .W36(W36TO84), .W37(W37TO84), .W38(W38TO84), .W39(W39TO84), .W40(W40TO84), .W41(W41TO84), .W42(W42TO84), .W43(W43TO84), .W44(W44TO84), .W45(W45TO84), .W46(W46TO84), .W47(W47TO84), .W48(W48TO84), .W49(W49TO84), .W50(W50TO84), .W51(W51TO84), .W52(W52TO84), .W53(W53TO84), .W54(W54TO84), .W55(W55TO84), .W56(W56TO84), .W57(W57TO84), .W58(W58TO84), .W59(W59TO84), .W60(W60TO84), .W61(W61TO84), .W62(W62TO84), .W63(W63TO84)) neuron84(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out84));
neuron64in #(.W0(W0TO85), .W1(W1TO85), .W2(W2TO85), .W3(W3TO85), .W4(W4TO85), .W5(W5TO85), .W6(W6TO85), .W7(W7TO85), .W8(W8TO85), .W9(W9TO85), .W10(W10TO85), .W11(W11TO85), .W12(W12TO85), .W13(W13TO85), .W14(W14TO85), .W15(W15TO85), .W16(W16TO85), .W17(W17TO85), .W18(W18TO85), .W19(W19TO85), .W20(W20TO85), .W21(W21TO85), .W22(W22TO85), .W23(W23TO85), .W24(W24TO85), .W25(W25TO85), .W26(W26TO85), .W27(W27TO85), .W28(W28TO85), .W29(W29TO85), .W30(W30TO85), .W31(W31TO85), .W32(W32TO85), .W33(W33TO85), .W34(W34TO85), .W35(W35TO85), .W36(W36TO85), .W37(W37TO85), .W38(W38TO85), .W39(W39TO85), .W40(W40TO85), .W41(W41TO85), .W42(W42TO85), .W43(W43TO85), .W44(W44TO85), .W45(W45TO85), .W46(W46TO85), .W47(W47TO85), .W48(W48TO85), .W49(W49TO85), .W50(W50TO85), .W51(W51TO85), .W52(W52TO85), .W53(W53TO85), .W54(W54TO85), .W55(W55TO85), .W56(W56TO85), .W57(W57TO85), .W58(W58TO85), .W59(W59TO85), .W60(W60TO85), .W61(W61TO85), .W62(W62TO85), .W63(W63TO85)) neuron85(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out85));
neuron64in #(.W0(W0TO86), .W1(W1TO86), .W2(W2TO86), .W3(W3TO86), .W4(W4TO86), .W5(W5TO86), .W6(W6TO86), .W7(W7TO86), .W8(W8TO86), .W9(W9TO86), .W10(W10TO86), .W11(W11TO86), .W12(W12TO86), .W13(W13TO86), .W14(W14TO86), .W15(W15TO86), .W16(W16TO86), .W17(W17TO86), .W18(W18TO86), .W19(W19TO86), .W20(W20TO86), .W21(W21TO86), .W22(W22TO86), .W23(W23TO86), .W24(W24TO86), .W25(W25TO86), .W26(W26TO86), .W27(W27TO86), .W28(W28TO86), .W29(W29TO86), .W30(W30TO86), .W31(W31TO86), .W32(W32TO86), .W33(W33TO86), .W34(W34TO86), .W35(W35TO86), .W36(W36TO86), .W37(W37TO86), .W38(W38TO86), .W39(W39TO86), .W40(W40TO86), .W41(W41TO86), .W42(W42TO86), .W43(W43TO86), .W44(W44TO86), .W45(W45TO86), .W46(W46TO86), .W47(W47TO86), .W48(W48TO86), .W49(W49TO86), .W50(W50TO86), .W51(W51TO86), .W52(W52TO86), .W53(W53TO86), .W54(W54TO86), .W55(W55TO86), .W56(W56TO86), .W57(W57TO86), .W58(W58TO86), .W59(W59TO86), .W60(W60TO86), .W61(W61TO86), .W62(W62TO86), .W63(W63TO86)) neuron86(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out86));
neuron64in #(.W0(W0TO87), .W1(W1TO87), .W2(W2TO87), .W3(W3TO87), .W4(W4TO87), .W5(W5TO87), .W6(W6TO87), .W7(W7TO87), .W8(W8TO87), .W9(W9TO87), .W10(W10TO87), .W11(W11TO87), .W12(W12TO87), .W13(W13TO87), .W14(W14TO87), .W15(W15TO87), .W16(W16TO87), .W17(W17TO87), .W18(W18TO87), .W19(W19TO87), .W20(W20TO87), .W21(W21TO87), .W22(W22TO87), .W23(W23TO87), .W24(W24TO87), .W25(W25TO87), .W26(W26TO87), .W27(W27TO87), .W28(W28TO87), .W29(W29TO87), .W30(W30TO87), .W31(W31TO87), .W32(W32TO87), .W33(W33TO87), .W34(W34TO87), .W35(W35TO87), .W36(W36TO87), .W37(W37TO87), .W38(W38TO87), .W39(W39TO87), .W40(W40TO87), .W41(W41TO87), .W42(W42TO87), .W43(W43TO87), .W44(W44TO87), .W45(W45TO87), .W46(W46TO87), .W47(W47TO87), .W48(W48TO87), .W49(W49TO87), .W50(W50TO87), .W51(W51TO87), .W52(W52TO87), .W53(W53TO87), .W54(W54TO87), .W55(W55TO87), .W56(W56TO87), .W57(W57TO87), .W58(W58TO87), .W59(W59TO87), .W60(W60TO87), .W61(W61TO87), .W62(W62TO87), .W63(W63TO87)) neuron87(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out87));
neuron64in #(.W0(W0TO88), .W1(W1TO88), .W2(W2TO88), .W3(W3TO88), .W4(W4TO88), .W5(W5TO88), .W6(W6TO88), .W7(W7TO88), .W8(W8TO88), .W9(W9TO88), .W10(W10TO88), .W11(W11TO88), .W12(W12TO88), .W13(W13TO88), .W14(W14TO88), .W15(W15TO88), .W16(W16TO88), .W17(W17TO88), .W18(W18TO88), .W19(W19TO88), .W20(W20TO88), .W21(W21TO88), .W22(W22TO88), .W23(W23TO88), .W24(W24TO88), .W25(W25TO88), .W26(W26TO88), .W27(W27TO88), .W28(W28TO88), .W29(W29TO88), .W30(W30TO88), .W31(W31TO88), .W32(W32TO88), .W33(W33TO88), .W34(W34TO88), .W35(W35TO88), .W36(W36TO88), .W37(W37TO88), .W38(W38TO88), .W39(W39TO88), .W40(W40TO88), .W41(W41TO88), .W42(W42TO88), .W43(W43TO88), .W44(W44TO88), .W45(W45TO88), .W46(W46TO88), .W47(W47TO88), .W48(W48TO88), .W49(W49TO88), .W50(W50TO88), .W51(W51TO88), .W52(W52TO88), .W53(W53TO88), .W54(W54TO88), .W55(W55TO88), .W56(W56TO88), .W57(W57TO88), .W58(W58TO88), .W59(W59TO88), .W60(W60TO88), .W61(W61TO88), .W62(W62TO88), .W63(W63TO88)) neuron88(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out88));
neuron64in #(.W0(W0TO89), .W1(W1TO89), .W2(W2TO89), .W3(W3TO89), .W4(W4TO89), .W5(W5TO89), .W6(W6TO89), .W7(W7TO89), .W8(W8TO89), .W9(W9TO89), .W10(W10TO89), .W11(W11TO89), .W12(W12TO89), .W13(W13TO89), .W14(W14TO89), .W15(W15TO89), .W16(W16TO89), .W17(W17TO89), .W18(W18TO89), .W19(W19TO89), .W20(W20TO89), .W21(W21TO89), .W22(W22TO89), .W23(W23TO89), .W24(W24TO89), .W25(W25TO89), .W26(W26TO89), .W27(W27TO89), .W28(W28TO89), .W29(W29TO89), .W30(W30TO89), .W31(W31TO89), .W32(W32TO89), .W33(W33TO89), .W34(W34TO89), .W35(W35TO89), .W36(W36TO89), .W37(W37TO89), .W38(W38TO89), .W39(W39TO89), .W40(W40TO89), .W41(W41TO89), .W42(W42TO89), .W43(W43TO89), .W44(W44TO89), .W45(W45TO89), .W46(W46TO89), .W47(W47TO89), .W48(W48TO89), .W49(W49TO89), .W50(W50TO89), .W51(W51TO89), .W52(W52TO89), .W53(W53TO89), .W54(W54TO89), .W55(W55TO89), .W56(W56TO89), .W57(W57TO89), .W58(W58TO89), .W59(W59TO89), .W60(W60TO89), .W61(W61TO89), .W62(W62TO89), .W63(W63TO89)) neuron89(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out89));
neuron64in #(.W0(W0TO90), .W1(W1TO90), .W2(W2TO90), .W3(W3TO90), .W4(W4TO90), .W5(W5TO90), .W6(W6TO90), .W7(W7TO90), .W8(W8TO90), .W9(W9TO90), .W10(W10TO90), .W11(W11TO90), .W12(W12TO90), .W13(W13TO90), .W14(W14TO90), .W15(W15TO90), .W16(W16TO90), .W17(W17TO90), .W18(W18TO90), .W19(W19TO90), .W20(W20TO90), .W21(W21TO90), .W22(W22TO90), .W23(W23TO90), .W24(W24TO90), .W25(W25TO90), .W26(W26TO90), .W27(W27TO90), .W28(W28TO90), .W29(W29TO90), .W30(W30TO90), .W31(W31TO90), .W32(W32TO90), .W33(W33TO90), .W34(W34TO90), .W35(W35TO90), .W36(W36TO90), .W37(W37TO90), .W38(W38TO90), .W39(W39TO90), .W40(W40TO90), .W41(W41TO90), .W42(W42TO90), .W43(W43TO90), .W44(W44TO90), .W45(W45TO90), .W46(W46TO90), .W47(W47TO90), .W48(W48TO90), .W49(W49TO90), .W50(W50TO90), .W51(W51TO90), .W52(W52TO90), .W53(W53TO90), .W54(W54TO90), .W55(W55TO90), .W56(W56TO90), .W57(W57TO90), .W58(W58TO90), .W59(W59TO90), .W60(W60TO90), .W61(W61TO90), .W62(W62TO90), .W63(W63TO90)) neuron90(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out90));
neuron64in #(.W0(W0TO91), .W1(W1TO91), .W2(W2TO91), .W3(W3TO91), .W4(W4TO91), .W5(W5TO91), .W6(W6TO91), .W7(W7TO91), .W8(W8TO91), .W9(W9TO91), .W10(W10TO91), .W11(W11TO91), .W12(W12TO91), .W13(W13TO91), .W14(W14TO91), .W15(W15TO91), .W16(W16TO91), .W17(W17TO91), .W18(W18TO91), .W19(W19TO91), .W20(W20TO91), .W21(W21TO91), .W22(W22TO91), .W23(W23TO91), .W24(W24TO91), .W25(W25TO91), .W26(W26TO91), .W27(W27TO91), .W28(W28TO91), .W29(W29TO91), .W30(W30TO91), .W31(W31TO91), .W32(W32TO91), .W33(W33TO91), .W34(W34TO91), .W35(W35TO91), .W36(W36TO91), .W37(W37TO91), .W38(W38TO91), .W39(W39TO91), .W40(W40TO91), .W41(W41TO91), .W42(W42TO91), .W43(W43TO91), .W44(W44TO91), .W45(W45TO91), .W46(W46TO91), .W47(W47TO91), .W48(W48TO91), .W49(W49TO91), .W50(W50TO91), .W51(W51TO91), .W52(W52TO91), .W53(W53TO91), .W54(W54TO91), .W55(W55TO91), .W56(W56TO91), .W57(W57TO91), .W58(W58TO91), .W59(W59TO91), .W60(W60TO91), .W61(W61TO91), .W62(W62TO91), .W63(W63TO91)) neuron91(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out91));
neuron64in #(.W0(W0TO92), .W1(W1TO92), .W2(W2TO92), .W3(W3TO92), .W4(W4TO92), .W5(W5TO92), .W6(W6TO92), .W7(W7TO92), .W8(W8TO92), .W9(W9TO92), .W10(W10TO92), .W11(W11TO92), .W12(W12TO92), .W13(W13TO92), .W14(W14TO92), .W15(W15TO92), .W16(W16TO92), .W17(W17TO92), .W18(W18TO92), .W19(W19TO92), .W20(W20TO92), .W21(W21TO92), .W22(W22TO92), .W23(W23TO92), .W24(W24TO92), .W25(W25TO92), .W26(W26TO92), .W27(W27TO92), .W28(W28TO92), .W29(W29TO92), .W30(W30TO92), .W31(W31TO92), .W32(W32TO92), .W33(W33TO92), .W34(W34TO92), .W35(W35TO92), .W36(W36TO92), .W37(W37TO92), .W38(W38TO92), .W39(W39TO92), .W40(W40TO92), .W41(W41TO92), .W42(W42TO92), .W43(W43TO92), .W44(W44TO92), .W45(W45TO92), .W46(W46TO92), .W47(W47TO92), .W48(W48TO92), .W49(W49TO92), .W50(W50TO92), .W51(W51TO92), .W52(W52TO92), .W53(W53TO92), .W54(W54TO92), .W55(W55TO92), .W56(W56TO92), .W57(W57TO92), .W58(W58TO92), .W59(W59TO92), .W60(W60TO92), .W61(W61TO92), .W62(W62TO92), .W63(W63TO92)) neuron92(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out92));
neuron64in #(.W0(W0TO93), .W1(W1TO93), .W2(W2TO93), .W3(W3TO93), .W4(W4TO93), .W5(W5TO93), .W6(W6TO93), .W7(W7TO93), .W8(W8TO93), .W9(W9TO93), .W10(W10TO93), .W11(W11TO93), .W12(W12TO93), .W13(W13TO93), .W14(W14TO93), .W15(W15TO93), .W16(W16TO93), .W17(W17TO93), .W18(W18TO93), .W19(W19TO93), .W20(W20TO93), .W21(W21TO93), .W22(W22TO93), .W23(W23TO93), .W24(W24TO93), .W25(W25TO93), .W26(W26TO93), .W27(W27TO93), .W28(W28TO93), .W29(W29TO93), .W30(W30TO93), .W31(W31TO93), .W32(W32TO93), .W33(W33TO93), .W34(W34TO93), .W35(W35TO93), .W36(W36TO93), .W37(W37TO93), .W38(W38TO93), .W39(W39TO93), .W40(W40TO93), .W41(W41TO93), .W42(W42TO93), .W43(W43TO93), .W44(W44TO93), .W45(W45TO93), .W46(W46TO93), .W47(W47TO93), .W48(W48TO93), .W49(W49TO93), .W50(W50TO93), .W51(W51TO93), .W52(W52TO93), .W53(W53TO93), .W54(W54TO93), .W55(W55TO93), .W56(W56TO93), .W57(W57TO93), .W58(W58TO93), .W59(W59TO93), .W60(W60TO93), .W61(W61TO93), .W62(W62TO93), .W63(W63TO93)) neuron93(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out93));
neuron64in #(.W0(W0TO94), .W1(W1TO94), .W2(W2TO94), .W3(W3TO94), .W4(W4TO94), .W5(W5TO94), .W6(W6TO94), .W7(W7TO94), .W8(W8TO94), .W9(W9TO94), .W10(W10TO94), .W11(W11TO94), .W12(W12TO94), .W13(W13TO94), .W14(W14TO94), .W15(W15TO94), .W16(W16TO94), .W17(W17TO94), .W18(W18TO94), .W19(W19TO94), .W20(W20TO94), .W21(W21TO94), .W22(W22TO94), .W23(W23TO94), .W24(W24TO94), .W25(W25TO94), .W26(W26TO94), .W27(W27TO94), .W28(W28TO94), .W29(W29TO94), .W30(W30TO94), .W31(W31TO94), .W32(W32TO94), .W33(W33TO94), .W34(W34TO94), .W35(W35TO94), .W36(W36TO94), .W37(W37TO94), .W38(W38TO94), .W39(W39TO94), .W40(W40TO94), .W41(W41TO94), .W42(W42TO94), .W43(W43TO94), .W44(W44TO94), .W45(W45TO94), .W46(W46TO94), .W47(W47TO94), .W48(W48TO94), .W49(W49TO94), .W50(W50TO94), .W51(W51TO94), .W52(W52TO94), .W53(W53TO94), .W54(W54TO94), .W55(W55TO94), .W56(W56TO94), .W57(W57TO94), .W58(W58TO94), .W59(W59TO94), .W60(W60TO94), .W61(W61TO94), .W62(W62TO94), .W63(W63TO94)) neuron94(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out94));
neuron64in #(.W0(W0TO95), .W1(W1TO95), .W2(W2TO95), .W3(W3TO95), .W4(W4TO95), .W5(W5TO95), .W6(W6TO95), .W7(W7TO95), .W8(W8TO95), .W9(W9TO95), .W10(W10TO95), .W11(W11TO95), .W12(W12TO95), .W13(W13TO95), .W14(W14TO95), .W15(W15TO95), .W16(W16TO95), .W17(W17TO95), .W18(W18TO95), .W19(W19TO95), .W20(W20TO95), .W21(W21TO95), .W22(W22TO95), .W23(W23TO95), .W24(W24TO95), .W25(W25TO95), .W26(W26TO95), .W27(W27TO95), .W28(W28TO95), .W29(W29TO95), .W30(W30TO95), .W31(W31TO95), .W32(W32TO95), .W33(W33TO95), .W34(W34TO95), .W35(W35TO95), .W36(W36TO95), .W37(W37TO95), .W38(W38TO95), .W39(W39TO95), .W40(W40TO95), .W41(W41TO95), .W42(W42TO95), .W43(W43TO95), .W44(W44TO95), .W45(W45TO95), .W46(W46TO95), .W47(W47TO95), .W48(W48TO95), .W49(W49TO95), .W50(W50TO95), .W51(W51TO95), .W52(W52TO95), .W53(W53TO95), .W54(W54TO95), .W55(W55TO95), .W56(W56TO95), .W57(W57TO95), .W58(W58TO95), .W59(W59TO95), .W60(W60TO95), .W61(W61TO95), .W62(W62TO95), .W63(W63TO95)) neuron95(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out95));
neuron64in #(.W0(W0TO96), .W1(W1TO96), .W2(W2TO96), .W3(W3TO96), .W4(W4TO96), .W5(W5TO96), .W6(W6TO96), .W7(W7TO96), .W8(W8TO96), .W9(W9TO96), .W10(W10TO96), .W11(W11TO96), .W12(W12TO96), .W13(W13TO96), .W14(W14TO96), .W15(W15TO96), .W16(W16TO96), .W17(W17TO96), .W18(W18TO96), .W19(W19TO96), .W20(W20TO96), .W21(W21TO96), .W22(W22TO96), .W23(W23TO96), .W24(W24TO96), .W25(W25TO96), .W26(W26TO96), .W27(W27TO96), .W28(W28TO96), .W29(W29TO96), .W30(W30TO96), .W31(W31TO96), .W32(W32TO96), .W33(W33TO96), .W34(W34TO96), .W35(W35TO96), .W36(W36TO96), .W37(W37TO96), .W38(W38TO96), .W39(W39TO96), .W40(W40TO96), .W41(W41TO96), .W42(W42TO96), .W43(W43TO96), .W44(W44TO96), .W45(W45TO96), .W46(W46TO96), .W47(W47TO96), .W48(W48TO96), .W49(W49TO96), .W50(W50TO96), .W51(W51TO96), .W52(W52TO96), .W53(W53TO96), .W54(W54TO96), .W55(W55TO96), .W56(W56TO96), .W57(W57TO96), .W58(W58TO96), .W59(W59TO96), .W60(W60TO96), .W61(W61TO96), .W62(W62TO96), .W63(W63TO96)) neuron96(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out96));
neuron64in #(.W0(W0TO97), .W1(W1TO97), .W2(W2TO97), .W3(W3TO97), .W4(W4TO97), .W5(W5TO97), .W6(W6TO97), .W7(W7TO97), .W8(W8TO97), .W9(W9TO97), .W10(W10TO97), .W11(W11TO97), .W12(W12TO97), .W13(W13TO97), .W14(W14TO97), .W15(W15TO97), .W16(W16TO97), .W17(W17TO97), .W18(W18TO97), .W19(W19TO97), .W20(W20TO97), .W21(W21TO97), .W22(W22TO97), .W23(W23TO97), .W24(W24TO97), .W25(W25TO97), .W26(W26TO97), .W27(W27TO97), .W28(W28TO97), .W29(W29TO97), .W30(W30TO97), .W31(W31TO97), .W32(W32TO97), .W33(W33TO97), .W34(W34TO97), .W35(W35TO97), .W36(W36TO97), .W37(W37TO97), .W38(W38TO97), .W39(W39TO97), .W40(W40TO97), .W41(W41TO97), .W42(W42TO97), .W43(W43TO97), .W44(W44TO97), .W45(W45TO97), .W46(W46TO97), .W47(W47TO97), .W48(W48TO97), .W49(W49TO97), .W50(W50TO97), .W51(W51TO97), .W52(W52TO97), .W53(W53TO97), .W54(W54TO97), .W55(W55TO97), .W56(W56TO97), .W57(W57TO97), .W58(W58TO97), .W59(W59TO97), .W60(W60TO97), .W61(W61TO97), .W62(W62TO97), .W63(W63TO97)) neuron97(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out97));
neuron64in #(.W0(W0TO98), .W1(W1TO98), .W2(W2TO98), .W3(W3TO98), .W4(W4TO98), .W5(W5TO98), .W6(W6TO98), .W7(W7TO98), .W8(W8TO98), .W9(W9TO98), .W10(W10TO98), .W11(W11TO98), .W12(W12TO98), .W13(W13TO98), .W14(W14TO98), .W15(W15TO98), .W16(W16TO98), .W17(W17TO98), .W18(W18TO98), .W19(W19TO98), .W20(W20TO98), .W21(W21TO98), .W22(W22TO98), .W23(W23TO98), .W24(W24TO98), .W25(W25TO98), .W26(W26TO98), .W27(W27TO98), .W28(W28TO98), .W29(W29TO98), .W30(W30TO98), .W31(W31TO98), .W32(W32TO98), .W33(W33TO98), .W34(W34TO98), .W35(W35TO98), .W36(W36TO98), .W37(W37TO98), .W38(W38TO98), .W39(W39TO98), .W40(W40TO98), .W41(W41TO98), .W42(W42TO98), .W43(W43TO98), .W44(W44TO98), .W45(W45TO98), .W46(W46TO98), .W47(W47TO98), .W48(W48TO98), .W49(W49TO98), .W50(W50TO98), .W51(W51TO98), .W52(W52TO98), .W53(W53TO98), .W54(W54TO98), .W55(W55TO98), .W56(W56TO98), .W57(W57TO98), .W58(W58TO98), .W59(W59TO98), .W60(W60TO98), .W61(W61TO98), .W62(W62TO98), .W63(W63TO98)) neuron98(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out98));
neuron64in #(.W0(W0TO99), .W1(W1TO99), .W2(W2TO99), .W3(W3TO99), .W4(W4TO99), .W5(W5TO99), .W6(W6TO99), .W7(W7TO99), .W8(W8TO99), .W9(W9TO99), .W10(W10TO99), .W11(W11TO99), .W12(W12TO99), .W13(W13TO99), .W14(W14TO99), .W15(W15TO99), .W16(W16TO99), .W17(W17TO99), .W18(W18TO99), .W19(W19TO99), .W20(W20TO99), .W21(W21TO99), .W22(W22TO99), .W23(W23TO99), .W24(W24TO99), .W25(W25TO99), .W26(W26TO99), .W27(W27TO99), .W28(W28TO99), .W29(W29TO99), .W30(W30TO99), .W31(W31TO99), .W32(W32TO99), .W33(W33TO99), .W34(W34TO99), .W35(W35TO99), .W36(W36TO99), .W37(W37TO99), .W38(W38TO99), .W39(W39TO99), .W40(W40TO99), .W41(W41TO99), .W42(W42TO99), .W43(W43TO99), .W44(W44TO99), .W45(W45TO99), .W46(W46TO99), .W47(W47TO99), .W48(W48TO99), .W49(W49TO99), .W50(W50TO99), .W51(W51TO99), .W52(W52TO99), .W53(W53TO99), .W54(W54TO99), .W55(W55TO99), .W56(W56TO99), .W57(W57TO99), .W58(W58TO99), .W59(W59TO99), .W60(W60TO99), .W61(W61TO99), .W62(W62TO99), .W63(W63TO99)) neuron99(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out99));

endmodule

module layer100in10out(clk, rst, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, in65, in66, in67, in68, in69, in70, in71, in72, in73, in74, in75, in76, in77, in78, in79, in80, in81, in82, in83, in84, in85, in86, in87, in88, in89, in90, in91, in92, in93, in94, in95, in96, in97, in98, in99, out0, out1, out2, out3, out4, out5, out6, out7, out8, out9);

parameter W0TO0 = 0;
parameter W0TO1 = 0;
parameter W0TO2 = 0;
parameter W0TO3 = 0;
parameter W0TO4 = 0;
parameter W0TO5 = 0;
parameter W0TO6 = 0;
parameter W0TO7 = 0;
parameter W0TO8 = 0;
parameter W0TO9 = 0;
parameter W1TO0 = 0;
parameter W1TO1 = 0;
parameter W1TO2 = 0;
parameter W1TO3 = 0;
parameter W1TO4 = 0;
parameter W1TO5 = 0;
parameter W1TO6 = 0;
parameter W1TO7 = 0;
parameter W1TO8 = 0;
parameter W1TO9 = 0;
parameter W2TO0 = 0;
parameter W2TO1 = 0;
parameter W2TO2 = 0;
parameter W2TO3 = 0;
parameter W2TO4 = 0;
parameter W2TO5 = 0;
parameter W2TO6 = 0;
parameter W2TO7 = 0;
parameter W2TO8 = 0;
parameter W2TO9 = 0;
parameter W3TO0 = 0;
parameter W3TO1 = 0;
parameter W3TO2 = 0;
parameter W3TO3 = 0;
parameter W3TO4 = 0;
parameter W3TO5 = 0;
parameter W3TO6 = 0;
parameter W3TO7 = 0;
parameter W3TO8 = 0;
parameter W3TO9 = 0;
parameter W4TO0 = 0;
parameter W4TO1 = 0;
parameter W4TO2 = 0;
parameter W4TO3 = 0;
parameter W4TO4 = 0;
parameter W4TO5 = 0;
parameter W4TO6 = 0;
parameter W4TO7 = 0;
parameter W4TO8 = 0;
parameter W4TO9 = 0;
parameter W5TO0 = 0;
parameter W5TO1 = 0;
parameter W5TO2 = 0;
parameter W5TO3 = 0;
parameter W5TO4 = 0;
parameter W5TO5 = 0;
parameter W5TO6 = 0;
parameter W5TO7 = 0;
parameter W5TO8 = 0;
parameter W5TO9 = 0;
parameter W6TO0 = 0;
parameter W6TO1 = 0;
parameter W6TO2 = 0;
parameter W6TO3 = 0;
parameter W6TO4 = 0;
parameter W6TO5 = 0;
parameter W6TO6 = 0;
parameter W6TO7 = 0;
parameter W6TO8 = 0;
parameter W6TO9 = 0;
parameter W7TO0 = 0;
parameter W7TO1 = 0;
parameter W7TO2 = 0;
parameter W7TO3 = 0;
parameter W7TO4 = 0;
parameter W7TO5 = 0;
parameter W7TO6 = 0;
parameter W7TO7 = 0;
parameter W7TO8 = 0;
parameter W7TO9 = 0;
parameter W8TO0 = 0;
parameter W8TO1 = 0;
parameter W8TO2 = 0;
parameter W8TO3 = 0;
parameter W8TO4 = 0;
parameter W8TO5 = 0;
parameter W8TO6 = 0;
parameter W8TO7 = 0;
parameter W8TO8 = 0;
parameter W8TO9 = 0;
parameter W9TO0 = 0;
parameter W9TO1 = 0;
parameter W9TO2 = 0;
parameter W9TO3 = 0;
parameter W9TO4 = 0;
parameter W9TO5 = 0;
parameter W9TO6 = 0;
parameter W9TO7 = 0;
parameter W9TO8 = 0;
parameter W9TO9 = 0;
parameter W10TO0 = 0;
parameter W10TO1 = 0;
parameter W10TO2 = 0;
parameter W10TO3 = 0;
parameter W10TO4 = 0;
parameter W10TO5 = 0;
parameter W10TO6 = 0;
parameter W10TO7 = 0;
parameter W10TO8 = 0;
parameter W10TO9 = 0;
parameter W11TO0 = 0;
parameter W11TO1 = 0;
parameter W11TO2 = 0;
parameter W11TO3 = 0;
parameter W11TO4 = 0;
parameter W11TO5 = 0;
parameter W11TO6 = 0;
parameter W11TO7 = 0;
parameter W11TO8 = 0;
parameter W11TO9 = 0;
parameter W12TO0 = 0;
parameter W12TO1 = 0;
parameter W12TO2 = 0;
parameter W12TO3 = 0;
parameter W12TO4 = 0;
parameter W12TO5 = 0;
parameter W12TO6 = 0;
parameter W12TO7 = 0;
parameter W12TO8 = 0;
parameter W12TO9 = 0;
parameter W13TO0 = 0;
parameter W13TO1 = 0;
parameter W13TO2 = 0;
parameter W13TO3 = 0;
parameter W13TO4 = 0;
parameter W13TO5 = 0;
parameter W13TO6 = 0;
parameter W13TO7 = 0;
parameter W13TO8 = 0;
parameter W13TO9 = 0;
parameter W14TO0 = 0;
parameter W14TO1 = 0;
parameter W14TO2 = 0;
parameter W14TO3 = 0;
parameter W14TO4 = 0;
parameter W14TO5 = 0;
parameter W14TO6 = 0;
parameter W14TO7 = 0;
parameter W14TO8 = 0;
parameter W14TO9 = 0;
parameter W15TO0 = 0;
parameter W15TO1 = 0;
parameter W15TO2 = 0;
parameter W15TO3 = 0;
parameter W15TO4 = 0;
parameter W15TO5 = 0;
parameter W15TO6 = 0;
parameter W15TO7 = 0;
parameter W15TO8 = 0;
parameter W15TO9 = 0;
parameter W16TO0 = 0;
parameter W16TO1 = 0;
parameter W16TO2 = 0;
parameter W16TO3 = 0;
parameter W16TO4 = 0;
parameter W16TO5 = 0;
parameter W16TO6 = 0;
parameter W16TO7 = 0;
parameter W16TO8 = 0;
parameter W16TO9 = 0;
parameter W17TO0 = 0;
parameter W17TO1 = 0;
parameter W17TO2 = 0;
parameter W17TO3 = 0;
parameter W17TO4 = 0;
parameter W17TO5 = 0;
parameter W17TO6 = 0;
parameter W17TO7 = 0;
parameter W17TO8 = 0;
parameter W17TO9 = 0;
parameter W18TO0 = 0;
parameter W18TO1 = 0;
parameter W18TO2 = 0;
parameter W18TO3 = 0;
parameter W18TO4 = 0;
parameter W18TO5 = 0;
parameter W18TO6 = 0;
parameter W18TO7 = 0;
parameter W18TO8 = 0;
parameter W18TO9 = 0;
parameter W19TO0 = 0;
parameter W19TO1 = 0;
parameter W19TO2 = 0;
parameter W19TO3 = 0;
parameter W19TO4 = 0;
parameter W19TO5 = 0;
parameter W19TO6 = 0;
parameter W19TO7 = 0;
parameter W19TO8 = 0;
parameter W19TO9 = 0;
parameter W20TO0 = 0;
parameter W20TO1 = 0;
parameter W20TO2 = 0;
parameter W20TO3 = 0;
parameter W20TO4 = 0;
parameter W20TO5 = 0;
parameter W20TO6 = 0;
parameter W20TO7 = 0;
parameter W20TO8 = 0;
parameter W20TO9 = 0;
parameter W21TO0 = 0;
parameter W21TO1 = 0;
parameter W21TO2 = 0;
parameter W21TO3 = 0;
parameter W21TO4 = 0;
parameter W21TO5 = 0;
parameter W21TO6 = 0;
parameter W21TO7 = 0;
parameter W21TO8 = 0;
parameter W21TO9 = 0;
parameter W22TO0 = 0;
parameter W22TO1 = 0;
parameter W22TO2 = 0;
parameter W22TO3 = 0;
parameter W22TO4 = 0;
parameter W22TO5 = 0;
parameter W22TO6 = 0;
parameter W22TO7 = 0;
parameter W22TO8 = 0;
parameter W22TO9 = 0;
parameter W23TO0 = 0;
parameter W23TO1 = 0;
parameter W23TO2 = 0;
parameter W23TO3 = 0;
parameter W23TO4 = 0;
parameter W23TO5 = 0;
parameter W23TO6 = 0;
parameter W23TO7 = 0;
parameter W23TO8 = 0;
parameter W23TO9 = 0;
parameter W24TO0 = 0;
parameter W24TO1 = 0;
parameter W24TO2 = 0;
parameter W24TO3 = 0;
parameter W24TO4 = 0;
parameter W24TO5 = 0;
parameter W24TO6 = 0;
parameter W24TO7 = 0;
parameter W24TO8 = 0;
parameter W24TO9 = 0;
parameter W25TO0 = 0;
parameter W25TO1 = 0;
parameter W25TO2 = 0;
parameter W25TO3 = 0;
parameter W25TO4 = 0;
parameter W25TO5 = 0;
parameter W25TO6 = 0;
parameter W25TO7 = 0;
parameter W25TO8 = 0;
parameter W25TO9 = 0;
parameter W26TO0 = 0;
parameter W26TO1 = 0;
parameter W26TO2 = 0;
parameter W26TO3 = 0;
parameter W26TO4 = 0;
parameter W26TO5 = 0;
parameter W26TO6 = 0;
parameter W26TO7 = 0;
parameter W26TO8 = 0;
parameter W26TO9 = 0;
parameter W27TO0 = 0;
parameter W27TO1 = 0;
parameter W27TO2 = 0;
parameter W27TO3 = 0;
parameter W27TO4 = 0;
parameter W27TO5 = 0;
parameter W27TO6 = 0;
parameter W27TO7 = 0;
parameter W27TO8 = 0;
parameter W27TO9 = 0;
parameter W28TO0 = 0;
parameter W28TO1 = 0;
parameter W28TO2 = 0;
parameter W28TO3 = 0;
parameter W28TO4 = 0;
parameter W28TO5 = 0;
parameter W28TO6 = 0;
parameter W28TO7 = 0;
parameter W28TO8 = 0;
parameter W28TO9 = 0;
parameter W29TO0 = 0;
parameter W29TO1 = 0;
parameter W29TO2 = 0;
parameter W29TO3 = 0;
parameter W29TO4 = 0;
parameter W29TO5 = 0;
parameter W29TO6 = 0;
parameter W29TO7 = 0;
parameter W29TO8 = 0;
parameter W29TO9 = 0;
parameter W30TO0 = 0;
parameter W30TO1 = 0;
parameter W30TO2 = 0;
parameter W30TO3 = 0;
parameter W30TO4 = 0;
parameter W30TO5 = 0;
parameter W30TO6 = 0;
parameter W30TO7 = 0;
parameter W30TO8 = 0;
parameter W30TO9 = 0;
parameter W31TO0 = 0;
parameter W31TO1 = 0;
parameter W31TO2 = 0;
parameter W31TO3 = 0;
parameter W31TO4 = 0;
parameter W31TO5 = 0;
parameter W31TO6 = 0;
parameter W31TO7 = 0;
parameter W31TO8 = 0;
parameter W31TO9 = 0;
parameter W32TO0 = 0;
parameter W32TO1 = 0;
parameter W32TO2 = 0;
parameter W32TO3 = 0;
parameter W32TO4 = 0;
parameter W32TO5 = 0;
parameter W32TO6 = 0;
parameter W32TO7 = 0;
parameter W32TO8 = 0;
parameter W32TO9 = 0;
parameter W33TO0 = 0;
parameter W33TO1 = 0;
parameter W33TO2 = 0;
parameter W33TO3 = 0;
parameter W33TO4 = 0;
parameter W33TO5 = 0;
parameter W33TO6 = 0;
parameter W33TO7 = 0;
parameter W33TO8 = 0;
parameter W33TO9 = 0;
parameter W34TO0 = 0;
parameter W34TO1 = 0;
parameter W34TO2 = 0;
parameter W34TO3 = 0;
parameter W34TO4 = 0;
parameter W34TO5 = 0;
parameter W34TO6 = 0;
parameter W34TO7 = 0;
parameter W34TO8 = 0;
parameter W34TO9 = 0;
parameter W35TO0 = 0;
parameter W35TO1 = 0;
parameter W35TO2 = 0;
parameter W35TO3 = 0;
parameter W35TO4 = 0;
parameter W35TO5 = 0;
parameter W35TO6 = 0;
parameter W35TO7 = 0;
parameter W35TO8 = 0;
parameter W35TO9 = 0;
parameter W36TO0 = 0;
parameter W36TO1 = 0;
parameter W36TO2 = 0;
parameter W36TO3 = 0;
parameter W36TO4 = 0;
parameter W36TO5 = 0;
parameter W36TO6 = 0;
parameter W36TO7 = 0;
parameter W36TO8 = 0;
parameter W36TO9 = 0;
parameter W37TO0 = 0;
parameter W37TO1 = 0;
parameter W37TO2 = 0;
parameter W37TO3 = 0;
parameter W37TO4 = 0;
parameter W37TO5 = 0;
parameter W37TO6 = 0;
parameter W37TO7 = 0;
parameter W37TO8 = 0;
parameter W37TO9 = 0;
parameter W38TO0 = 0;
parameter W38TO1 = 0;
parameter W38TO2 = 0;
parameter W38TO3 = 0;
parameter W38TO4 = 0;
parameter W38TO5 = 0;
parameter W38TO6 = 0;
parameter W38TO7 = 0;
parameter W38TO8 = 0;
parameter W38TO9 = 0;
parameter W39TO0 = 0;
parameter W39TO1 = 0;
parameter W39TO2 = 0;
parameter W39TO3 = 0;
parameter W39TO4 = 0;
parameter W39TO5 = 0;
parameter W39TO6 = 0;
parameter W39TO7 = 0;
parameter W39TO8 = 0;
parameter W39TO9 = 0;
parameter W40TO0 = 0;
parameter W40TO1 = 0;
parameter W40TO2 = 0;
parameter W40TO3 = 0;
parameter W40TO4 = 0;
parameter W40TO5 = 0;
parameter W40TO6 = 0;
parameter W40TO7 = 0;
parameter W40TO8 = 0;
parameter W40TO9 = 0;
parameter W41TO0 = 0;
parameter W41TO1 = 0;
parameter W41TO2 = 0;
parameter W41TO3 = 0;
parameter W41TO4 = 0;
parameter W41TO5 = 0;
parameter W41TO6 = 0;
parameter W41TO7 = 0;
parameter W41TO8 = 0;
parameter W41TO9 = 0;
parameter W42TO0 = 0;
parameter W42TO1 = 0;
parameter W42TO2 = 0;
parameter W42TO3 = 0;
parameter W42TO4 = 0;
parameter W42TO5 = 0;
parameter W42TO6 = 0;
parameter W42TO7 = 0;
parameter W42TO8 = 0;
parameter W42TO9 = 0;
parameter W43TO0 = 0;
parameter W43TO1 = 0;
parameter W43TO2 = 0;
parameter W43TO3 = 0;
parameter W43TO4 = 0;
parameter W43TO5 = 0;
parameter W43TO6 = 0;
parameter W43TO7 = 0;
parameter W43TO8 = 0;
parameter W43TO9 = 0;
parameter W44TO0 = 0;
parameter W44TO1 = 0;
parameter W44TO2 = 0;
parameter W44TO3 = 0;
parameter W44TO4 = 0;
parameter W44TO5 = 0;
parameter W44TO6 = 0;
parameter W44TO7 = 0;
parameter W44TO8 = 0;
parameter W44TO9 = 0;
parameter W45TO0 = 0;
parameter W45TO1 = 0;
parameter W45TO2 = 0;
parameter W45TO3 = 0;
parameter W45TO4 = 0;
parameter W45TO5 = 0;
parameter W45TO6 = 0;
parameter W45TO7 = 0;
parameter W45TO8 = 0;
parameter W45TO9 = 0;
parameter W46TO0 = 0;
parameter W46TO1 = 0;
parameter W46TO2 = 0;
parameter W46TO3 = 0;
parameter W46TO4 = 0;
parameter W46TO5 = 0;
parameter W46TO6 = 0;
parameter W46TO7 = 0;
parameter W46TO8 = 0;
parameter W46TO9 = 0;
parameter W47TO0 = 0;
parameter W47TO1 = 0;
parameter W47TO2 = 0;
parameter W47TO3 = 0;
parameter W47TO4 = 0;
parameter W47TO5 = 0;
parameter W47TO6 = 0;
parameter W47TO7 = 0;
parameter W47TO8 = 0;
parameter W47TO9 = 0;
parameter W48TO0 = 0;
parameter W48TO1 = 0;
parameter W48TO2 = 0;
parameter W48TO3 = 0;
parameter W48TO4 = 0;
parameter W48TO5 = 0;
parameter W48TO6 = 0;
parameter W48TO7 = 0;
parameter W48TO8 = 0;
parameter W48TO9 = 0;
parameter W49TO0 = 0;
parameter W49TO1 = 0;
parameter W49TO2 = 0;
parameter W49TO3 = 0;
parameter W49TO4 = 0;
parameter W49TO5 = 0;
parameter W49TO6 = 0;
parameter W49TO7 = 0;
parameter W49TO8 = 0;
parameter W49TO9 = 0;
parameter W50TO0 = 0;
parameter W50TO1 = 0;
parameter W50TO2 = 0;
parameter W50TO3 = 0;
parameter W50TO4 = 0;
parameter W50TO5 = 0;
parameter W50TO6 = 0;
parameter W50TO7 = 0;
parameter W50TO8 = 0;
parameter W50TO9 = 0;
parameter W51TO0 = 0;
parameter W51TO1 = 0;
parameter W51TO2 = 0;
parameter W51TO3 = 0;
parameter W51TO4 = 0;
parameter W51TO5 = 0;
parameter W51TO6 = 0;
parameter W51TO7 = 0;
parameter W51TO8 = 0;
parameter W51TO9 = 0;
parameter W52TO0 = 0;
parameter W52TO1 = 0;
parameter W52TO2 = 0;
parameter W52TO3 = 0;
parameter W52TO4 = 0;
parameter W52TO5 = 0;
parameter W52TO6 = 0;
parameter W52TO7 = 0;
parameter W52TO8 = 0;
parameter W52TO9 = 0;
parameter W53TO0 = 0;
parameter W53TO1 = 0;
parameter W53TO2 = 0;
parameter W53TO3 = 0;
parameter W53TO4 = 0;
parameter W53TO5 = 0;
parameter W53TO6 = 0;
parameter W53TO7 = 0;
parameter W53TO8 = 0;
parameter W53TO9 = 0;
parameter W54TO0 = 0;
parameter W54TO1 = 0;
parameter W54TO2 = 0;
parameter W54TO3 = 0;
parameter W54TO4 = 0;
parameter W54TO5 = 0;
parameter W54TO6 = 0;
parameter W54TO7 = 0;
parameter W54TO8 = 0;
parameter W54TO9 = 0;
parameter W55TO0 = 0;
parameter W55TO1 = 0;
parameter W55TO2 = 0;
parameter W55TO3 = 0;
parameter W55TO4 = 0;
parameter W55TO5 = 0;
parameter W55TO6 = 0;
parameter W55TO7 = 0;
parameter W55TO8 = 0;
parameter W55TO9 = 0;
parameter W56TO0 = 0;
parameter W56TO1 = 0;
parameter W56TO2 = 0;
parameter W56TO3 = 0;
parameter W56TO4 = 0;
parameter W56TO5 = 0;
parameter W56TO6 = 0;
parameter W56TO7 = 0;
parameter W56TO8 = 0;
parameter W56TO9 = 0;
parameter W57TO0 = 0;
parameter W57TO1 = 0;
parameter W57TO2 = 0;
parameter W57TO3 = 0;
parameter W57TO4 = 0;
parameter W57TO5 = 0;
parameter W57TO6 = 0;
parameter W57TO7 = 0;
parameter W57TO8 = 0;
parameter W57TO9 = 0;
parameter W58TO0 = 0;
parameter W58TO1 = 0;
parameter W58TO2 = 0;
parameter W58TO3 = 0;
parameter W58TO4 = 0;
parameter W58TO5 = 0;
parameter W58TO6 = 0;
parameter W58TO7 = 0;
parameter W58TO8 = 0;
parameter W58TO9 = 0;
parameter W59TO0 = 0;
parameter W59TO1 = 0;
parameter W59TO2 = 0;
parameter W59TO3 = 0;
parameter W59TO4 = 0;
parameter W59TO5 = 0;
parameter W59TO6 = 0;
parameter W59TO7 = 0;
parameter W59TO8 = 0;
parameter W59TO9 = 0;
parameter W60TO0 = 0;
parameter W60TO1 = 0;
parameter W60TO2 = 0;
parameter W60TO3 = 0;
parameter W60TO4 = 0;
parameter W60TO5 = 0;
parameter W60TO6 = 0;
parameter W60TO7 = 0;
parameter W60TO8 = 0;
parameter W60TO9 = 0;
parameter W61TO0 = 0;
parameter W61TO1 = 0;
parameter W61TO2 = 0;
parameter W61TO3 = 0;
parameter W61TO4 = 0;
parameter W61TO5 = 0;
parameter W61TO6 = 0;
parameter W61TO7 = 0;
parameter W61TO8 = 0;
parameter W61TO9 = 0;
parameter W62TO0 = 0;
parameter W62TO1 = 0;
parameter W62TO2 = 0;
parameter W62TO3 = 0;
parameter W62TO4 = 0;
parameter W62TO5 = 0;
parameter W62TO6 = 0;
parameter W62TO7 = 0;
parameter W62TO8 = 0;
parameter W62TO9 = 0;
parameter W63TO0 = 0;
parameter W63TO1 = 0;
parameter W63TO2 = 0;
parameter W63TO3 = 0;
parameter W63TO4 = 0;
parameter W63TO5 = 0;
parameter W63TO6 = 0;
parameter W63TO7 = 0;
parameter W63TO8 = 0;
parameter W63TO9 = 0;
parameter W64TO0 = 0;
parameter W64TO1 = 0;
parameter W64TO2 = 0;
parameter W64TO3 = 0;
parameter W64TO4 = 0;
parameter W64TO5 = 0;
parameter W64TO6 = 0;
parameter W64TO7 = 0;
parameter W64TO8 = 0;
parameter W64TO9 = 0;
parameter W65TO0 = 0;
parameter W65TO1 = 0;
parameter W65TO2 = 0;
parameter W65TO3 = 0;
parameter W65TO4 = 0;
parameter W65TO5 = 0;
parameter W65TO6 = 0;
parameter W65TO7 = 0;
parameter W65TO8 = 0;
parameter W65TO9 = 0;
parameter W66TO0 = 0;
parameter W66TO1 = 0;
parameter W66TO2 = 0;
parameter W66TO3 = 0;
parameter W66TO4 = 0;
parameter W66TO5 = 0;
parameter W66TO6 = 0;
parameter W66TO7 = 0;
parameter W66TO8 = 0;
parameter W66TO9 = 0;
parameter W67TO0 = 0;
parameter W67TO1 = 0;
parameter W67TO2 = 0;
parameter W67TO3 = 0;
parameter W67TO4 = 0;
parameter W67TO5 = 0;
parameter W67TO6 = 0;
parameter W67TO7 = 0;
parameter W67TO8 = 0;
parameter W67TO9 = 0;
parameter W68TO0 = 0;
parameter W68TO1 = 0;
parameter W68TO2 = 0;
parameter W68TO3 = 0;
parameter W68TO4 = 0;
parameter W68TO5 = 0;
parameter W68TO6 = 0;
parameter W68TO7 = 0;
parameter W68TO8 = 0;
parameter W68TO9 = 0;
parameter W69TO0 = 0;
parameter W69TO1 = 0;
parameter W69TO2 = 0;
parameter W69TO3 = 0;
parameter W69TO4 = 0;
parameter W69TO5 = 0;
parameter W69TO6 = 0;
parameter W69TO7 = 0;
parameter W69TO8 = 0;
parameter W69TO9 = 0;
parameter W70TO0 = 0;
parameter W70TO1 = 0;
parameter W70TO2 = 0;
parameter W70TO3 = 0;
parameter W70TO4 = 0;
parameter W70TO5 = 0;
parameter W70TO6 = 0;
parameter W70TO7 = 0;
parameter W70TO8 = 0;
parameter W70TO9 = 0;
parameter W71TO0 = 0;
parameter W71TO1 = 0;
parameter W71TO2 = 0;
parameter W71TO3 = 0;
parameter W71TO4 = 0;
parameter W71TO5 = 0;
parameter W71TO6 = 0;
parameter W71TO7 = 0;
parameter W71TO8 = 0;
parameter W71TO9 = 0;
parameter W72TO0 = 0;
parameter W72TO1 = 0;
parameter W72TO2 = 0;
parameter W72TO3 = 0;
parameter W72TO4 = 0;
parameter W72TO5 = 0;
parameter W72TO6 = 0;
parameter W72TO7 = 0;
parameter W72TO8 = 0;
parameter W72TO9 = 0;
parameter W73TO0 = 0;
parameter W73TO1 = 0;
parameter W73TO2 = 0;
parameter W73TO3 = 0;
parameter W73TO4 = 0;
parameter W73TO5 = 0;
parameter W73TO6 = 0;
parameter W73TO7 = 0;
parameter W73TO8 = 0;
parameter W73TO9 = 0;
parameter W74TO0 = 0;
parameter W74TO1 = 0;
parameter W74TO2 = 0;
parameter W74TO3 = 0;
parameter W74TO4 = 0;
parameter W74TO5 = 0;
parameter W74TO6 = 0;
parameter W74TO7 = 0;
parameter W74TO8 = 0;
parameter W74TO9 = 0;
parameter W75TO0 = 0;
parameter W75TO1 = 0;
parameter W75TO2 = 0;
parameter W75TO3 = 0;
parameter W75TO4 = 0;
parameter W75TO5 = 0;
parameter W75TO6 = 0;
parameter W75TO7 = 0;
parameter W75TO8 = 0;
parameter W75TO9 = 0;
parameter W76TO0 = 0;
parameter W76TO1 = 0;
parameter W76TO2 = 0;
parameter W76TO3 = 0;
parameter W76TO4 = 0;
parameter W76TO5 = 0;
parameter W76TO6 = 0;
parameter W76TO7 = 0;
parameter W76TO8 = 0;
parameter W76TO9 = 0;
parameter W77TO0 = 0;
parameter W77TO1 = 0;
parameter W77TO2 = 0;
parameter W77TO3 = 0;
parameter W77TO4 = 0;
parameter W77TO5 = 0;
parameter W77TO6 = 0;
parameter W77TO7 = 0;
parameter W77TO8 = 0;
parameter W77TO9 = 0;
parameter W78TO0 = 0;
parameter W78TO1 = 0;
parameter W78TO2 = 0;
parameter W78TO3 = 0;
parameter W78TO4 = 0;
parameter W78TO5 = 0;
parameter W78TO6 = 0;
parameter W78TO7 = 0;
parameter W78TO8 = 0;
parameter W78TO9 = 0;
parameter W79TO0 = 0;
parameter W79TO1 = 0;
parameter W79TO2 = 0;
parameter W79TO3 = 0;
parameter W79TO4 = 0;
parameter W79TO5 = 0;
parameter W79TO6 = 0;
parameter W79TO7 = 0;
parameter W79TO8 = 0;
parameter W79TO9 = 0;
parameter W80TO0 = 0;
parameter W80TO1 = 0;
parameter W80TO2 = 0;
parameter W80TO3 = 0;
parameter W80TO4 = 0;
parameter W80TO5 = 0;
parameter W80TO6 = 0;
parameter W80TO7 = 0;
parameter W80TO8 = 0;
parameter W80TO9 = 0;
parameter W81TO0 = 0;
parameter W81TO1 = 0;
parameter W81TO2 = 0;
parameter W81TO3 = 0;
parameter W81TO4 = 0;
parameter W81TO5 = 0;
parameter W81TO6 = 0;
parameter W81TO7 = 0;
parameter W81TO8 = 0;
parameter W81TO9 = 0;
parameter W82TO0 = 0;
parameter W82TO1 = 0;
parameter W82TO2 = 0;
parameter W82TO3 = 0;
parameter W82TO4 = 0;
parameter W82TO5 = 0;
parameter W82TO6 = 0;
parameter W82TO7 = 0;
parameter W82TO8 = 0;
parameter W82TO9 = 0;
parameter W83TO0 = 0;
parameter W83TO1 = 0;
parameter W83TO2 = 0;
parameter W83TO3 = 0;
parameter W83TO4 = 0;
parameter W83TO5 = 0;
parameter W83TO6 = 0;
parameter W83TO7 = 0;
parameter W83TO8 = 0;
parameter W83TO9 = 0;
parameter W84TO0 = 0;
parameter W84TO1 = 0;
parameter W84TO2 = 0;
parameter W84TO3 = 0;
parameter W84TO4 = 0;
parameter W84TO5 = 0;
parameter W84TO6 = 0;
parameter W84TO7 = 0;
parameter W84TO8 = 0;
parameter W84TO9 = 0;
parameter W85TO0 = 0;
parameter W85TO1 = 0;
parameter W85TO2 = 0;
parameter W85TO3 = 0;
parameter W85TO4 = 0;
parameter W85TO5 = 0;
parameter W85TO6 = 0;
parameter W85TO7 = 0;
parameter W85TO8 = 0;
parameter W85TO9 = 0;
parameter W86TO0 = 0;
parameter W86TO1 = 0;
parameter W86TO2 = 0;
parameter W86TO3 = 0;
parameter W86TO4 = 0;
parameter W86TO5 = 0;
parameter W86TO6 = 0;
parameter W86TO7 = 0;
parameter W86TO8 = 0;
parameter W86TO9 = 0;
parameter W87TO0 = 0;
parameter W87TO1 = 0;
parameter W87TO2 = 0;
parameter W87TO3 = 0;
parameter W87TO4 = 0;
parameter W87TO5 = 0;
parameter W87TO6 = 0;
parameter W87TO7 = 0;
parameter W87TO8 = 0;
parameter W87TO9 = 0;
parameter W88TO0 = 0;
parameter W88TO1 = 0;
parameter W88TO2 = 0;
parameter W88TO3 = 0;
parameter W88TO4 = 0;
parameter W88TO5 = 0;
parameter W88TO6 = 0;
parameter W88TO7 = 0;
parameter W88TO8 = 0;
parameter W88TO9 = 0;
parameter W89TO0 = 0;
parameter W89TO1 = 0;
parameter W89TO2 = 0;
parameter W89TO3 = 0;
parameter W89TO4 = 0;
parameter W89TO5 = 0;
parameter W89TO6 = 0;
parameter W89TO7 = 0;
parameter W89TO8 = 0;
parameter W89TO9 = 0;
parameter W90TO0 = 0;
parameter W90TO1 = 0;
parameter W90TO2 = 0;
parameter W90TO3 = 0;
parameter W90TO4 = 0;
parameter W90TO5 = 0;
parameter W90TO6 = 0;
parameter W90TO7 = 0;
parameter W90TO8 = 0;
parameter W90TO9 = 0;
parameter W91TO0 = 0;
parameter W91TO1 = 0;
parameter W91TO2 = 0;
parameter W91TO3 = 0;
parameter W91TO4 = 0;
parameter W91TO5 = 0;
parameter W91TO6 = 0;
parameter W91TO7 = 0;
parameter W91TO8 = 0;
parameter W91TO9 = 0;
parameter W92TO0 = 0;
parameter W92TO1 = 0;
parameter W92TO2 = 0;
parameter W92TO3 = 0;
parameter W92TO4 = 0;
parameter W92TO5 = 0;
parameter W92TO6 = 0;
parameter W92TO7 = 0;
parameter W92TO8 = 0;
parameter W92TO9 = 0;
parameter W93TO0 = 0;
parameter W93TO1 = 0;
parameter W93TO2 = 0;
parameter W93TO3 = 0;
parameter W93TO4 = 0;
parameter W93TO5 = 0;
parameter W93TO6 = 0;
parameter W93TO7 = 0;
parameter W93TO8 = 0;
parameter W93TO9 = 0;
parameter W94TO0 = 0;
parameter W94TO1 = 0;
parameter W94TO2 = 0;
parameter W94TO3 = 0;
parameter W94TO4 = 0;
parameter W94TO5 = 0;
parameter W94TO6 = 0;
parameter W94TO7 = 0;
parameter W94TO8 = 0;
parameter W94TO9 = 0;
parameter W95TO0 = 0;
parameter W95TO1 = 0;
parameter W95TO2 = 0;
parameter W95TO3 = 0;
parameter W95TO4 = 0;
parameter W95TO5 = 0;
parameter W95TO6 = 0;
parameter W95TO7 = 0;
parameter W95TO8 = 0;
parameter W95TO9 = 0;
parameter W96TO0 = 0;
parameter W96TO1 = 0;
parameter W96TO2 = 0;
parameter W96TO3 = 0;
parameter W96TO4 = 0;
parameter W96TO5 = 0;
parameter W96TO6 = 0;
parameter W96TO7 = 0;
parameter W96TO8 = 0;
parameter W96TO9 = 0;
parameter W97TO0 = 0;
parameter W97TO1 = 0;
parameter W97TO2 = 0;
parameter W97TO3 = 0;
parameter W97TO4 = 0;
parameter W97TO5 = 0;
parameter W97TO6 = 0;
parameter W97TO7 = 0;
parameter W97TO8 = 0;
parameter W97TO9 = 0;
parameter W98TO0 = 0;
parameter W98TO1 = 0;
parameter W98TO2 = 0;
parameter W98TO3 = 0;
parameter W98TO4 = 0;
parameter W98TO5 = 0;
parameter W98TO6 = 0;
parameter W98TO7 = 0;
parameter W98TO8 = 0;
parameter W98TO9 = 0;
parameter W99TO0 = 0;
parameter W99TO1 = 0;
parameter W99TO2 = 0;
parameter W99TO3 = 0;
parameter W99TO4 = 0;
parameter W99TO5 = 0;
parameter W99TO6 = 0;
parameter W99TO7 = 0;
parameter W99TO8 = 0;
parameter W99TO9 = 0;

input wire clk;
input wire rst;

input signed [15:0] in0;
input signed [15:0] in1;
input signed [15:0] in2;
input signed [15:0] in3;
input signed [15:0] in4;
input signed [15:0] in5;
input signed [15:0] in6;
input signed [15:0] in7;
input signed [15:0] in8;
input signed [15:0] in9;
input signed [15:0] in10;
input signed [15:0] in11;
input signed [15:0] in12;
input signed [15:0] in13;
input signed [15:0] in14;
input signed [15:0] in15;
input signed [15:0] in16;
input signed [15:0] in17;
input signed [15:0] in18;
input signed [15:0] in19;
input signed [15:0] in20;
input signed [15:0] in21;
input signed [15:0] in22;
input signed [15:0] in23;
input signed [15:0] in24;
input signed [15:0] in25;
input signed [15:0] in26;
input signed [15:0] in27;
input signed [15:0] in28;
input signed [15:0] in29;
input signed [15:0] in30;
input signed [15:0] in31;
input signed [15:0] in32;
input signed [15:0] in33;
input signed [15:0] in34;
input signed [15:0] in35;
input signed [15:0] in36;
input signed [15:0] in37;
input signed [15:0] in38;
input signed [15:0] in39;
input signed [15:0] in40;
input signed [15:0] in41;
input signed [15:0] in42;
input signed [15:0] in43;
input signed [15:0] in44;
input signed [15:0] in45;
input signed [15:0] in46;
input signed [15:0] in47;
input signed [15:0] in48;
input signed [15:0] in49;
input signed [15:0] in50;
input signed [15:0] in51;
input signed [15:0] in52;
input signed [15:0] in53;
input signed [15:0] in54;
input signed [15:0] in55;
input signed [15:0] in56;
input signed [15:0] in57;
input signed [15:0] in58;
input signed [15:0] in59;
input signed [15:0] in60;
input signed [15:0] in61;
input signed [15:0] in62;
input signed [15:0] in63;
input signed [15:0] in64;
input signed [15:0] in65;
input signed [15:0] in66;
input signed [15:0] in67;
input signed [15:0] in68;
input signed [15:0] in69;
input signed [15:0] in70;
input signed [15:0] in71;
input signed [15:0] in72;
input signed [15:0] in73;
input signed [15:0] in74;
input signed [15:0] in75;
input signed [15:0] in76;
input signed [15:0] in77;
input signed [15:0] in78;
input signed [15:0] in79;
input signed [15:0] in80;
input signed [15:0] in81;
input signed [15:0] in82;
input signed [15:0] in83;
input signed [15:0] in84;
input signed [15:0] in85;
input signed [15:0] in86;
input signed [15:0] in87;
input signed [15:0] in88;
input signed [15:0] in89;
input signed [15:0] in90;
input signed [15:0] in91;
input signed [15:0] in92;
input signed [15:0] in93;
input signed [15:0] in94;
input signed [15:0] in95;
input signed [15:0] in96;
input signed [15:0] in97;
input signed [15:0] in98;
input signed [15:0] in99;

output signed [15:0] out0;
output signed [15:0] out1;
output signed [15:0] out2;
output signed [15:0] out3;
output signed [15:0] out4;
output signed [15:0] out5;
output signed [15:0] out6;
output signed [15:0] out7;
output signed [15:0] out8;
output signed [15:0] out9;

neuron100in #(.W0(W0TO0), .W1(W1TO0), .W2(W2TO0), .W3(W3TO0), .W4(W4TO0), .W5(W5TO0), .W6(W6TO0), .W7(W7TO0), .W8(W8TO0), .W9(W9TO0), .W10(W10TO0), .W11(W11TO0), .W12(W12TO0), .W13(W13TO0), .W14(W14TO0), .W15(W15TO0), .W16(W16TO0), .W17(W17TO0), .W18(W18TO0), .W19(W19TO0), .W20(W20TO0), .W21(W21TO0), .W22(W22TO0), .W23(W23TO0), .W24(W24TO0), .W25(W25TO0), .W26(W26TO0), .W27(W27TO0), .W28(W28TO0), .W29(W29TO0), .W30(W30TO0), .W31(W31TO0), .W32(W32TO0), .W33(W33TO0), .W34(W34TO0), .W35(W35TO0), .W36(W36TO0), .W37(W37TO0), .W38(W38TO0), .W39(W39TO0), .W40(W40TO0), .W41(W41TO0), .W42(W42TO0), .W43(W43TO0), .W44(W44TO0), .W45(W45TO0), .W46(W46TO0), .W47(W47TO0), .W48(W48TO0), .W49(W49TO0), .W50(W50TO0), .W51(W51TO0), .W52(W52TO0), .W53(W53TO0), .W54(W54TO0), .W55(W55TO0), .W56(W56TO0), .W57(W57TO0), .W58(W58TO0), .W59(W59TO0), .W60(W60TO0), .W61(W61TO0), .W62(W62TO0), .W63(W63TO0), .W64(W64TO0), .W65(W65TO0), .W66(W66TO0), .W67(W67TO0), .W68(W68TO0), .W69(W69TO0), .W70(W70TO0), .W71(W71TO0), .W72(W72TO0), .W73(W73TO0), .W74(W74TO0), .W75(W75TO0), .W76(W76TO0), .W77(W77TO0), .W78(W78TO0), .W79(W79TO0), .W80(W80TO0), .W81(W81TO0), .W82(W82TO0), .W83(W83TO0), .W84(W84TO0), .W85(W85TO0), .W86(W86TO0), .W87(W87TO0), .W88(W88TO0), .W89(W89TO0), .W90(W90TO0), .W91(W91TO0), .W92(W92TO0), .W93(W93TO0), .W94(W94TO0), .W95(W95TO0), .W96(W96TO0), .W97(W97TO0), .W98(W98TO0), .W99(W99TO0)) neuron0(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .in65(in65), .in66(in66), .in67(in67), .in68(in68), .in69(in69), .in70(in70), .in71(in71), .in72(in72), .in73(in73), .in74(in74), .in75(in75), .in76(in76), .in77(in77), .in78(in78), .in79(in79), .in80(in80), .in81(in81), .in82(in82), .in83(in83), .in84(in84), .in85(in85), .in86(in86), .in87(in87), .in88(in88), .in89(in89), .in90(in90), .in91(in91), .in92(in92), .in93(in93), .in94(in94), .in95(in95), .in96(in96), .in97(in97), .in98(in98), .in99(in99), .out(out0));
neuron100in #(.W0(W0TO1), .W1(W1TO1), .W2(W2TO1), .W3(W3TO1), .W4(W4TO1), .W5(W5TO1), .W6(W6TO1), .W7(W7TO1), .W8(W8TO1), .W9(W9TO1), .W10(W10TO1), .W11(W11TO1), .W12(W12TO1), .W13(W13TO1), .W14(W14TO1), .W15(W15TO1), .W16(W16TO1), .W17(W17TO1), .W18(W18TO1), .W19(W19TO1), .W20(W20TO1), .W21(W21TO1), .W22(W22TO1), .W23(W23TO1), .W24(W24TO1), .W25(W25TO1), .W26(W26TO1), .W27(W27TO1), .W28(W28TO1), .W29(W29TO1), .W30(W30TO1), .W31(W31TO1), .W32(W32TO1), .W33(W33TO1), .W34(W34TO1), .W35(W35TO1), .W36(W36TO1), .W37(W37TO1), .W38(W38TO1), .W39(W39TO1), .W40(W40TO1), .W41(W41TO1), .W42(W42TO1), .W43(W43TO1), .W44(W44TO1), .W45(W45TO1), .W46(W46TO1), .W47(W47TO1), .W48(W48TO1), .W49(W49TO1), .W50(W50TO1), .W51(W51TO1), .W52(W52TO1), .W53(W53TO1), .W54(W54TO1), .W55(W55TO1), .W56(W56TO1), .W57(W57TO1), .W58(W58TO1), .W59(W59TO1), .W60(W60TO1), .W61(W61TO1), .W62(W62TO1), .W63(W63TO1), .W64(W64TO1), .W65(W65TO1), .W66(W66TO1), .W67(W67TO1), .W68(W68TO1), .W69(W69TO1), .W70(W70TO1), .W71(W71TO1), .W72(W72TO1), .W73(W73TO1), .W74(W74TO1), .W75(W75TO1), .W76(W76TO1), .W77(W77TO1), .W78(W78TO1), .W79(W79TO1), .W80(W80TO1), .W81(W81TO1), .W82(W82TO1), .W83(W83TO1), .W84(W84TO1), .W85(W85TO1), .W86(W86TO1), .W87(W87TO1), .W88(W88TO1), .W89(W89TO1), .W90(W90TO1), .W91(W91TO1), .W92(W92TO1), .W93(W93TO1), .W94(W94TO1), .W95(W95TO1), .W96(W96TO1), .W97(W97TO1), .W98(W98TO1), .W99(W99TO1)) neuron1(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .in65(in65), .in66(in66), .in67(in67), .in68(in68), .in69(in69), .in70(in70), .in71(in71), .in72(in72), .in73(in73), .in74(in74), .in75(in75), .in76(in76), .in77(in77), .in78(in78), .in79(in79), .in80(in80), .in81(in81), .in82(in82), .in83(in83), .in84(in84), .in85(in85), .in86(in86), .in87(in87), .in88(in88), .in89(in89), .in90(in90), .in91(in91), .in92(in92), .in93(in93), .in94(in94), .in95(in95), .in96(in96), .in97(in97), .in98(in98), .in99(in99), .out(out1));
neuron100in #(.W0(W0TO2), .W1(W1TO2), .W2(W2TO2), .W3(W3TO2), .W4(W4TO2), .W5(W5TO2), .W6(W6TO2), .W7(W7TO2), .W8(W8TO2), .W9(W9TO2), .W10(W10TO2), .W11(W11TO2), .W12(W12TO2), .W13(W13TO2), .W14(W14TO2), .W15(W15TO2), .W16(W16TO2), .W17(W17TO2), .W18(W18TO2), .W19(W19TO2), .W20(W20TO2), .W21(W21TO2), .W22(W22TO2), .W23(W23TO2), .W24(W24TO2), .W25(W25TO2), .W26(W26TO2), .W27(W27TO2), .W28(W28TO2), .W29(W29TO2), .W30(W30TO2), .W31(W31TO2), .W32(W32TO2), .W33(W33TO2), .W34(W34TO2), .W35(W35TO2), .W36(W36TO2), .W37(W37TO2), .W38(W38TO2), .W39(W39TO2), .W40(W40TO2), .W41(W41TO2), .W42(W42TO2), .W43(W43TO2), .W44(W44TO2), .W45(W45TO2), .W46(W46TO2), .W47(W47TO2), .W48(W48TO2), .W49(W49TO2), .W50(W50TO2), .W51(W51TO2), .W52(W52TO2), .W53(W53TO2), .W54(W54TO2), .W55(W55TO2), .W56(W56TO2), .W57(W57TO2), .W58(W58TO2), .W59(W59TO2), .W60(W60TO2), .W61(W61TO2), .W62(W62TO2), .W63(W63TO2), .W64(W64TO2), .W65(W65TO2), .W66(W66TO2), .W67(W67TO2), .W68(W68TO2), .W69(W69TO2), .W70(W70TO2), .W71(W71TO2), .W72(W72TO2), .W73(W73TO2), .W74(W74TO2), .W75(W75TO2), .W76(W76TO2), .W77(W77TO2), .W78(W78TO2), .W79(W79TO2), .W80(W80TO2), .W81(W81TO2), .W82(W82TO2), .W83(W83TO2), .W84(W84TO2), .W85(W85TO2), .W86(W86TO2), .W87(W87TO2), .W88(W88TO2), .W89(W89TO2), .W90(W90TO2), .W91(W91TO2), .W92(W92TO2), .W93(W93TO2), .W94(W94TO2), .W95(W95TO2), .W96(W96TO2), .W97(W97TO2), .W98(W98TO2), .W99(W99TO2)) neuron2(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .in65(in65), .in66(in66), .in67(in67), .in68(in68), .in69(in69), .in70(in70), .in71(in71), .in72(in72), .in73(in73), .in74(in74), .in75(in75), .in76(in76), .in77(in77), .in78(in78), .in79(in79), .in80(in80), .in81(in81), .in82(in82), .in83(in83), .in84(in84), .in85(in85), .in86(in86), .in87(in87), .in88(in88), .in89(in89), .in90(in90), .in91(in91), .in92(in92), .in93(in93), .in94(in94), .in95(in95), .in96(in96), .in97(in97), .in98(in98), .in99(in99), .out(out2));
neuron100in #(.W0(W0TO3), .W1(W1TO3), .W2(W2TO3), .W3(W3TO3), .W4(W4TO3), .W5(W5TO3), .W6(W6TO3), .W7(W7TO3), .W8(W8TO3), .W9(W9TO3), .W10(W10TO3), .W11(W11TO3), .W12(W12TO3), .W13(W13TO3), .W14(W14TO3), .W15(W15TO3), .W16(W16TO3), .W17(W17TO3), .W18(W18TO3), .W19(W19TO3), .W20(W20TO3), .W21(W21TO3), .W22(W22TO3), .W23(W23TO3), .W24(W24TO3), .W25(W25TO3), .W26(W26TO3), .W27(W27TO3), .W28(W28TO3), .W29(W29TO3), .W30(W30TO3), .W31(W31TO3), .W32(W32TO3), .W33(W33TO3), .W34(W34TO3), .W35(W35TO3), .W36(W36TO3), .W37(W37TO3), .W38(W38TO3), .W39(W39TO3), .W40(W40TO3), .W41(W41TO3), .W42(W42TO3), .W43(W43TO3), .W44(W44TO3), .W45(W45TO3), .W46(W46TO3), .W47(W47TO3), .W48(W48TO3), .W49(W49TO3), .W50(W50TO3), .W51(W51TO3), .W52(W52TO3), .W53(W53TO3), .W54(W54TO3), .W55(W55TO3), .W56(W56TO3), .W57(W57TO3), .W58(W58TO3), .W59(W59TO3), .W60(W60TO3), .W61(W61TO3), .W62(W62TO3), .W63(W63TO3), .W64(W64TO3), .W65(W65TO3), .W66(W66TO3), .W67(W67TO3), .W68(W68TO3), .W69(W69TO3), .W70(W70TO3), .W71(W71TO3), .W72(W72TO3), .W73(W73TO3), .W74(W74TO3), .W75(W75TO3), .W76(W76TO3), .W77(W77TO3), .W78(W78TO3), .W79(W79TO3), .W80(W80TO3), .W81(W81TO3), .W82(W82TO3), .W83(W83TO3), .W84(W84TO3), .W85(W85TO3), .W86(W86TO3), .W87(W87TO3), .W88(W88TO3), .W89(W89TO3), .W90(W90TO3), .W91(W91TO3), .W92(W92TO3), .W93(W93TO3), .W94(W94TO3), .W95(W95TO3), .W96(W96TO3), .W97(W97TO3), .W98(W98TO3), .W99(W99TO3)) neuron3(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .in65(in65), .in66(in66), .in67(in67), .in68(in68), .in69(in69), .in70(in70), .in71(in71), .in72(in72), .in73(in73), .in74(in74), .in75(in75), .in76(in76), .in77(in77), .in78(in78), .in79(in79), .in80(in80), .in81(in81), .in82(in82), .in83(in83), .in84(in84), .in85(in85), .in86(in86), .in87(in87), .in88(in88), .in89(in89), .in90(in90), .in91(in91), .in92(in92), .in93(in93), .in94(in94), .in95(in95), .in96(in96), .in97(in97), .in98(in98), .in99(in99), .out(out3));
neuron100in #(.W0(W0TO4), .W1(W1TO4), .W2(W2TO4), .W3(W3TO4), .W4(W4TO4), .W5(W5TO4), .W6(W6TO4), .W7(W7TO4), .W8(W8TO4), .W9(W9TO4), .W10(W10TO4), .W11(W11TO4), .W12(W12TO4), .W13(W13TO4), .W14(W14TO4), .W15(W15TO4), .W16(W16TO4), .W17(W17TO4), .W18(W18TO4), .W19(W19TO4), .W20(W20TO4), .W21(W21TO4), .W22(W22TO4), .W23(W23TO4), .W24(W24TO4), .W25(W25TO4), .W26(W26TO4), .W27(W27TO4), .W28(W28TO4), .W29(W29TO4), .W30(W30TO4), .W31(W31TO4), .W32(W32TO4), .W33(W33TO4), .W34(W34TO4), .W35(W35TO4), .W36(W36TO4), .W37(W37TO4), .W38(W38TO4), .W39(W39TO4), .W40(W40TO4), .W41(W41TO4), .W42(W42TO4), .W43(W43TO4), .W44(W44TO4), .W45(W45TO4), .W46(W46TO4), .W47(W47TO4), .W48(W48TO4), .W49(W49TO4), .W50(W50TO4), .W51(W51TO4), .W52(W52TO4), .W53(W53TO4), .W54(W54TO4), .W55(W55TO4), .W56(W56TO4), .W57(W57TO4), .W58(W58TO4), .W59(W59TO4), .W60(W60TO4), .W61(W61TO4), .W62(W62TO4), .W63(W63TO4), .W64(W64TO4), .W65(W65TO4), .W66(W66TO4), .W67(W67TO4), .W68(W68TO4), .W69(W69TO4), .W70(W70TO4), .W71(W71TO4), .W72(W72TO4), .W73(W73TO4), .W74(W74TO4), .W75(W75TO4), .W76(W76TO4), .W77(W77TO4), .W78(W78TO4), .W79(W79TO4), .W80(W80TO4), .W81(W81TO4), .W82(W82TO4), .W83(W83TO4), .W84(W84TO4), .W85(W85TO4), .W86(W86TO4), .W87(W87TO4), .W88(W88TO4), .W89(W89TO4), .W90(W90TO4), .W91(W91TO4), .W92(W92TO4), .W93(W93TO4), .W94(W94TO4), .W95(W95TO4), .W96(W96TO4), .W97(W97TO4), .W98(W98TO4), .W99(W99TO4)) neuron4(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .in65(in65), .in66(in66), .in67(in67), .in68(in68), .in69(in69), .in70(in70), .in71(in71), .in72(in72), .in73(in73), .in74(in74), .in75(in75), .in76(in76), .in77(in77), .in78(in78), .in79(in79), .in80(in80), .in81(in81), .in82(in82), .in83(in83), .in84(in84), .in85(in85), .in86(in86), .in87(in87), .in88(in88), .in89(in89), .in90(in90), .in91(in91), .in92(in92), .in93(in93), .in94(in94), .in95(in95), .in96(in96), .in97(in97), .in98(in98), .in99(in99), .out(out4));
neuron100in #(.W0(W0TO5), .W1(W1TO5), .W2(W2TO5), .W3(W3TO5), .W4(W4TO5), .W5(W5TO5), .W6(W6TO5), .W7(W7TO5), .W8(W8TO5), .W9(W9TO5), .W10(W10TO5), .W11(W11TO5), .W12(W12TO5), .W13(W13TO5), .W14(W14TO5), .W15(W15TO5), .W16(W16TO5), .W17(W17TO5), .W18(W18TO5), .W19(W19TO5), .W20(W20TO5), .W21(W21TO5), .W22(W22TO5), .W23(W23TO5), .W24(W24TO5), .W25(W25TO5), .W26(W26TO5), .W27(W27TO5), .W28(W28TO5), .W29(W29TO5), .W30(W30TO5), .W31(W31TO5), .W32(W32TO5), .W33(W33TO5), .W34(W34TO5), .W35(W35TO5), .W36(W36TO5), .W37(W37TO5), .W38(W38TO5), .W39(W39TO5), .W40(W40TO5), .W41(W41TO5), .W42(W42TO5), .W43(W43TO5), .W44(W44TO5), .W45(W45TO5), .W46(W46TO5), .W47(W47TO5), .W48(W48TO5), .W49(W49TO5), .W50(W50TO5), .W51(W51TO5), .W52(W52TO5), .W53(W53TO5), .W54(W54TO5), .W55(W55TO5), .W56(W56TO5), .W57(W57TO5), .W58(W58TO5), .W59(W59TO5), .W60(W60TO5), .W61(W61TO5), .W62(W62TO5), .W63(W63TO5), .W64(W64TO5), .W65(W65TO5), .W66(W66TO5), .W67(W67TO5), .W68(W68TO5), .W69(W69TO5), .W70(W70TO5), .W71(W71TO5), .W72(W72TO5), .W73(W73TO5), .W74(W74TO5), .W75(W75TO5), .W76(W76TO5), .W77(W77TO5), .W78(W78TO5), .W79(W79TO5), .W80(W80TO5), .W81(W81TO5), .W82(W82TO5), .W83(W83TO5), .W84(W84TO5), .W85(W85TO5), .W86(W86TO5), .W87(W87TO5), .W88(W88TO5), .W89(W89TO5), .W90(W90TO5), .W91(W91TO5), .W92(W92TO5), .W93(W93TO5), .W94(W94TO5), .W95(W95TO5), .W96(W96TO5), .W97(W97TO5), .W98(W98TO5), .W99(W99TO5)) neuron5(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .in65(in65), .in66(in66), .in67(in67), .in68(in68), .in69(in69), .in70(in70), .in71(in71), .in72(in72), .in73(in73), .in74(in74), .in75(in75), .in76(in76), .in77(in77), .in78(in78), .in79(in79), .in80(in80), .in81(in81), .in82(in82), .in83(in83), .in84(in84), .in85(in85), .in86(in86), .in87(in87), .in88(in88), .in89(in89), .in90(in90), .in91(in91), .in92(in92), .in93(in93), .in94(in94), .in95(in95), .in96(in96), .in97(in97), .in98(in98), .in99(in99), .out(out5));
neuron100in #(.W0(W0TO6), .W1(W1TO6), .W2(W2TO6), .W3(W3TO6), .W4(W4TO6), .W5(W5TO6), .W6(W6TO6), .W7(W7TO6), .W8(W8TO6), .W9(W9TO6), .W10(W10TO6), .W11(W11TO6), .W12(W12TO6), .W13(W13TO6), .W14(W14TO6), .W15(W15TO6), .W16(W16TO6), .W17(W17TO6), .W18(W18TO6), .W19(W19TO6), .W20(W20TO6), .W21(W21TO6), .W22(W22TO6), .W23(W23TO6), .W24(W24TO6), .W25(W25TO6), .W26(W26TO6), .W27(W27TO6), .W28(W28TO6), .W29(W29TO6), .W30(W30TO6), .W31(W31TO6), .W32(W32TO6), .W33(W33TO6), .W34(W34TO6), .W35(W35TO6), .W36(W36TO6), .W37(W37TO6), .W38(W38TO6), .W39(W39TO6), .W40(W40TO6), .W41(W41TO6), .W42(W42TO6), .W43(W43TO6), .W44(W44TO6), .W45(W45TO6), .W46(W46TO6), .W47(W47TO6), .W48(W48TO6), .W49(W49TO6), .W50(W50TO6), .W51(W51TO6), .W52(W52TO6), .W53(W53TO6), .W54(W54TO6), .W55(W55TO6), .W56(W56TO6), .W57(W57TO6), .W58(W58TO6), .W59(W59TO6), .W60(W60TO6), .W61(W61TO6), .W62(W62TO6), .W63(W63TO6), .W64(W64TO6), .W65(W65TO6), .W66(W66TO6), .W67(W67TO6), .W68(W68TO6), .W69(W69TO6), .W70(W70TO6), .W71(W71TO6), .W72(W72TO6), .W73(W73TO6), .W74(W74TO6), .W75(W75TO6), .W76(W76TO6), .W77(W77TO6), .W78(W78TO6), .W79(W79TO6), .W80(W80TO6), .W81(W81TO6), .W82(W82TO6), .W83(W83TO6), .W84(W84TO6), .W85(W85TO6), .W86(W86TO6), .W87(W87TO6), .W88(W88TO6), .W89(W89TO6), .W90(W90TO6), .W91(W91TO6), .W92(W92TO6), .W93(W93TO6), .W94(W94TO6), .W95(W95TO6), .W96(W96TO6), .W97(W97TO6), .W98(W98TO6), .W99(W99TO6)) neuron6(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .in65(in65), .in66(in66), .in67(in67), .in68(in68), .in69(in69), .in70(in70), .in71(in71), .in72(in72), .in73(in73), .in74(in74), .in75(in75), .in76(in76), .in77(in77), .in78(in78), .in79(in79), .in80(in80), .in81(in81), .in82(in82), .in83(in83), .in84(in84), .in85(in85), .in86(in86), .in87(in87), .in88(in88), .in89(in89), .in90(in90), .in91(in91), .in92(in92), .in93(in93), .in94(in94), .in95(in95), .in96(in96), .in97(in97), .in98(in98), .in99(in99), .out(out6));
neuron100in #(.W0(W0TO7), .W1(W1TO7), .W2(W2TO7), .W3(W3TO7), .W4(W4TO7), .W5(W5TO7), .W6(W6TO7), .W7(W7TO7), .W8(W8TO7), .W9(W9TO7), .W10(W10TO7), .W11(W11TO7), .W12(W12TO7), .W13(W13TO7), .W14(W14TO7), .W15(W15TO7), .W16(W16TO7), .W17(W17TO7), .W18(W18TO7), .W19(W19TO7), .W20(W20TO7), .W21(W21TO7), .W22(W22TO7), .W23(W23TO7), .W24(W24TO7), .W25(W25TO7), .W26(W26TO7), .W27(W27TO7), .W28(W28TO7), .W29(W29TO7), .W30(W30TO7), .W31(W31TO7), .W32(W32TO7), .W33(W33TO7), .W34(W34TO7), .W35(W35TO7), .W36(W36TO7), .W37(W37TO7), .W38(W38TO7), .W39(W39TO7), .W40(W40TO7), .W41(W41TO7), .W42(W42TO7), .W43(W43TO7), .W44(W44TO7), .W45(W45TO7), .W46(W46TO7), .W47(W47TO7), .W48(W48TO7), .W49(W49TO7), .W50(W50TO7), .W51(W51TO7), .W52(W52TO7), .W53(W53TO7), .W54(W54TO7), .W55(W55TO7), .W56(W56TO7), .W57(W57TO7), .W58(W58TO7), .W59(W59TO7), .W60(W60TO7), .W61(W61TO7), .W62(W62TO7), .W63(W63TO7), .W64(W64TO7), .W65(W65TO7), .W66(W66TO7), .W67(W67TO7), .W68(W68TO7), .W69(W69TO7), .W70(W70TO7), .W71(W71TO7), .W72(W72TO7), .W73(W73TO7), .W74(W74TO7), .W75(W75TO7), .W76(W76TO7), .W77(W77TO7), .W78(W78TO7), .W79(W79TO7), .W80(W80TO7), .W81(W81TO7), .W82(W82TO7), .W83(W83TO7), .W84(W84TO7), .W85(W85TO7), .W86(W86TO7), .W87(W87TO7), .W88(W88TO7), .W89(W89TO7), .W90(W90TO7), .W91(W91TO7), .W92(W92TO7), .W93(W93TO7), .W94(W94TO7), .W95(W95TO7), .W96(W96TO7), .W97(W97TO7), .W98(W98TO7), .W99(W99TO7)) neuron7(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .in65(in65), .in66(in66), .in67(in67), .in68(in68), .in69(in69), .in70(in70), .in71(in71), .in72(in72), .in73(in73), .in74(in74), .in75(in75), .in76(in76), .in77(in77), .in78(in78), .in79(in79), .in80(in80), .in81(in81), .in82(in82), .in83(in83), .in84(in84), .in85(in85), .in86(in86), .in87(in87), .in88(in88), .in89(in89), .in90(in90), .in91(in91), .in92(in92), .in93(in93), .in94(in94), .in95(in95), .in96(in96), .in97(in97), .in98(in98), .in99(in99), .out(out7));
neuron100in #(.W0(W0TO8), .W1(W1TO8), .W2(W2TO8), .W3(W3TO8), .W4(W4TO8), .W5(W5TO8), .W6(W6TO8), .W7(W7TO8), .W8(W8TO8), .W9(W9TO8), .W10(W10TO8), .W11(W11TO8), .W12(W12TO8), .W13(W13TO8), .W14(W14TO8), .W15(W15TO8), .W16(W16TO8), .W17(W17TO8), .W18(W18TO8), .W19(W19TO8), .W20(W20TO8), .W21(W21TO8), .W22(W22TO8), .W23(W23TO8), .W24(W24TO8), .W25(W25TO8), .W26(W26TO8), .W27(W27TO8), .W28(W28TO8), .W29(W29TO8), .W30(W30TO8), .W31(W31TO8), .W32(W32TO8), .W33(W33TO8), .W34(W34TO8), .W35(W35TO8), .W36(W36TO8), .W37(W37TO8), .W38(W38TO8), .W39(W39TO8), .W40(W40TO8), .W41(W41TO8), .W42(W42TO8), .W43(W43TO8), .W44(W44TO8), .W45(W45TO8), .W46(W46TO8), .W47(W47TO8), .W48(W48TO8), .W49(W49TO8), .W50(W50TO8), .W51(W51TO8), .W52(W52TO8), .W53(W53TO8), .W54(W54TO8), .W55(W55TO8), .W56(W56TO8), .W57(W57TO8), .W58(W58TO8), .W59(W59TO8), .W60(W60TO8), .W61(W61TO8), .W62(W62TO8), .W63(W63TO8), .W64(W64TO8), .W65(W65TO8), .W66(W66TO8), .W67(W67TO8), .W68(W68TO8), .W69(W69TO8), .W70(W70TO8), .W71(W71TO8), .W72(W72TO8), .W73(W73TO8), .W74(W74TO8), .W75(W75TO8), .W76(W76TO8), .W77(W77TO8), .W78(W78TO8), .W79(W79TO8), .W80(W80TO8), .W81(W81TO8), .W82(W82TO8), .W83(W83TO8), .W84(W84TO8), .W85(W85TO8), .W86(W86TO8), .W87(W87TO8), .W88(W88TO8), .W89(W89TO8), .W90(W90TO8), .W91(W91TO8), .W92(W92TO8), .W93(W93TO8), .W94(W94TO8), .W95(W95TO8), .W96(W96TO8), .W97(W97TO8), .W98(W98TO8), .W99(W99TO8)) neuron8(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .in65(in65), .in66(in66), .in67(in67), .in68(in68), .in69(in69), .in70(in70), .in71(in71), .in72(in72), .in73(in73), .in74(in74), .in75(in75), .in76(in76), .in77(in77), .in78(in78), .in79(in79), .in80(in80), .in81(in81), .in82(in82), .in83(in83), .in84(in84), .in85(in85), .in86(in86), .in87(in87), .in88(in88), .in89(in89), .in90(in90), .in91(in91), .in92(in92), .in93(in93), .in94(in94), .in95(in95), .in96(in96), .in97(in97), .in98(in98), .in99(in99), .out(out8));
neuron100in #(.W0(W0TO9), .W1(W1TO9), .W2(W2TO9), .W3(W3TO9), .W4(W4TO9), .W5(W5TO9), .W6(W6TO9), .W7(W7TO9), .W8(W8TO9), .W9(W9TO9), .W10(W10TO9), .W11(W11TO9), .W12(W12TO9), .W13(W13TO9), .W14(W14TO9), .W15(W15TO9), .W16(W16TO9), .W17(W17TO9), .W18(W18TO9), .W19(W19TO9), .W20(W20TO9), .W21(W21TO9), .W22(W22TO9), .W23(W23TO9), .W24(W24TO9), .W25(W25TO9), .W26(W26TO9), .W27(W27TO9), .W28(W28TO9), .W29(W29TO9), .W30(W30TO9), .W31(W31TO9), .W32(W32TO9), .W33(W33TO9), .W34(W34TO9), .W35(W35TO9), .W36(W36TO9), .W37(W37TO9), .W38(W38TO9), .W39(W39TO9), .W40(W40TO9), .W41(W41TO9), .W42(W42TO9), .W43(W43TO9), .W44(W44TO9), .W45(W45TO9), .W46(W46TO9), .W47(W47TO9), .W48(W48TO9), .W49(W49TO9), .W50(W50TO9), .W51(W51TO9), .W52(W52TO9), .W53(W53TO9), .W54(W54TO9), .W55(W55TO9), .W56(W56TO9), .W57(W57TO9), .W58(W58TO9), .W59(W59TO9), .W60(W60TO9), .W61(W61TO9), .W62(W62TO9), .W63(W63TO9), .W64(W64TO9), .W65(W65TO9), .W66(W66TO9), .W67(W67TO9), .W68(W68TO9), .W69(W69TO9), .W70(W70TO9), .W71(W71TO9), .W72(W72TO9), .W73(W73TO9), .W74(W74TO9), .W75(W75TO9), .W76(W76TO9), .W77(W77TO9), .W78(W78TO9), .W79(W79TO9), .W80(W80TO9), .W81(W81TO9), .W82(W82TO9), .W83(W83TO9), .W84(W84TO9), .W85(W85TO9), .W86(W86TO9), .W87(W87TO9), .W88(W88TO9), .W89(W89TO9), .W90(W90TO9), .W91(W91TO9), .W92(W92TO9), .W93(W93TO9), .W94(W94TO9), .W95(W95TO9), .W96(W96TO9), .W97(W97TO9), .W98(W98TO9), .W99(W99TO9)) neuron9(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .in65(in65), .in66(in66), .in67(in67), .in68(in68), .in69(in69), .in70(in70), .in71(in71), .in72(in72), .in73(in73), .in74(in74), .in75(in75), .in76(in76), .in77(in77), .in78(in78), .in79(in79), .in80(in80), .in81(in81), .in82(in82), .in83(in83), .in84(in84), .in85(in85), .in86(in86), .in87(in87), .in88(in88), .in89(in89), .in90(in90), .in91(in91), .in92(in92), .in93(in93), .in94(in94), .in95(in95), .in96(in96), .in97(in97), .in98(in98), .in99(in99), .out(out9));

endmodule

module network(clk, rst, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, out0, out1, out2, out3, out4, out5, out6, out7, out8, out9);

input wire clk;
input wire rst;

input signed [15:0] in0;
input signed [15:0] in1;
input signed [15:0] in2;
input signed [15:0] in3;
input signed [15:0] in4;
input signed [15:0] in5;
input signed [15:0] in6;
input signed [15:0] in7;
input signed [15:0] in8;
input signed [15:0] in9;
input signed [15:0] in10;
input signed [15:0] in11;
input signed [15:0] in12;
input signed [15:0] in13;
input signed [15:0] in14;
input signed [15:0] in15;
input signed [15:0] in16;
input signed [15:0] in17;
input signed [15:0] in18;
input signed [15:0] in19;
input signed [15:0] in20;
input signed [15:0] in21;
input signed [15:0] in22;
input signed [15:0] in23;
input signed [15:0] in24;
input signed [15:0] in25;
input signed [15:0] in26;
input signed [15:0] in27;
input signed [15:0] in28;
input signed [15:0] in29;
input signed [15:0] in30;
input signed [15:0] in31;
input signed [15:0] in32;
input signed [15:0] in33;
input signed [15:0] in34;
input signed [15:0] in35;
input signed [15:0] in36;
input signed [15:0] in37;
input signed [15:0] in38;
input signed [15:0] in39;
input signed [15:0] in40;
input signed [15:0] in41;
input signed [15:0] in42;
input signed [15:0] in43;
input signed [15:0] in44;
input signed [15:0] in45;
input signed [15:0] in46;
input signed [15:0] in47;
input signed [15:0] in48;
input signed [15:0] in49;
input signed [15:0] in50;
input signed [15:0] in51;
input signed [15:0] in52;
input signed [15:0] in53;
input signed [15:0] in54;
input signed [15:0] in55;
input signed [15:0] in56;
input signed [15:0] in57;
input signed [15:0] in58;
input signed [15:0] in59;
input signed [15:0] in60;
input signed [15:0] in61;
input signed [15:0] in62;
input signed [15:0] in63;

output signed [15:0] out0;
output signed [15:0] out1;
output signed [15:0] out2;
output signed [15:0] out3;
output signed [15:0] out4;
output signed [15:0] out5;
output signed [15:0] out6;
output signed [15:0] out7;
output signed [15:0] out8;
output signed [15:0] out9;

wire[15:0] con0[0:99];

layer64in100out #(.W0TO0(-145), .W0TO1(75), .W0TO2(114), .W0TO3(-22), .W0TO4(-127), .W0TO5(86), .W0TO6(-156), .W0TO7(146), .W0TO8(187), .W0TO9(-31), .W0TO10(53), .W0TO11(72), .W0TO12(-125), .W0TO13(-187), .W0TO14(-158), .W0TO15(-15), .W0TO16(167), .W0TO17(40), .W0TO18(-166), .W0TO19(-171), .W0TO20(66), .W0TO21(-183), .W0TO22(43), .W0TO23(-84), .W0TO24(102), .W0TO25(4), .W0TO26(24), .W0TO27(-170), .W0TO28(82), .W0TO29(8), .W0TO30(-95), .W0TO31(-152), .W0TO32(-45), .W0TO33(-177), .W0TO34(30), .W0TO35(95), .W0TO36(2), .W0TO37(-165), .W0TO38(-179), .W0TO39(47), .W0TO40(116), .W0TO41(-157), .W0TO42(20), .W0TO43(34), .W0TO44(-17), .W0TO45(23), .W0TO46(-73), .W0TO47(6), .W0TO48(-82), .W0TO49(140), .W0TO50(-146), .W0TO51(-148), .W0TO52(-113), .W0TO53(107), .W0TO54(29), .W0TO55(117), .W0TO56(74), .W0TO57(100), .W0TO58(86), .W0TO59(63), .W0TO60(-187), .W0TO61(30), .W0TO62(-47), .W0TO63(81), .W0TO64(33), .W0TO65(26), .W0TO66(90), .W0TO67(1), .W0TO68(120), .W0TO69(28), .W0TO70(-164), .W0TO71(138), .W0TO72(-189), .W0TO73(-86), .W0TO74(-106), .W0TO75(173), .W0TO76(81), .W0TO77(-53), .W0TO78(34), .W0TO79(100), .W0TO80(-91), .W0TO81(16), .W0TO82(-4), .W0TO83(-11), .W0TO84(-99), .W0TO85(20), .W0TO86(-112), .W0TO87(-42), .W0TO88(85), .W0TO89(96), .W0TO90(57), .W0TO91(-62), .W0TO92(-103), .W0TO93(-182), .W0TO94(113), .W0TO95(118), .W0TO96(118), .W0TO97(-140), .W0TO98(-88), .W0TO99(-57), .W1TO0(-155), .W1TO1(177), .W1TO2(87), .W1TO3(-164), .W1TO4(-187), .W1TO5(-172), .W1TO6(-18), .W1TO7(-150), .W1TO8(135), .W1TO9(-151), .W1TO10(90), .W1TO11(-171), .W1TO12(149), .W1TO13(-103), .W1TO14(-57), .W1TO15(13), .W1TO16(-41), .W1TO17(-153), .W1TO18(-69), .W1TO19(86), .W1TO20(-96), .W1TO21(162), .W1TO22(180), .W1TO23(-181), .W1TO24(29), .W1TO25(-124), .W1TO26(35), .W1TO27(130), .W1TO28(56), .W1TO29(52), .W1TO30(9), .W1TO31(-16), .W1TO32(-93), .W1TO33(98), .W1TO34(99), .W1TO35(102), .W1TO36(-198), .W1TO37(18), .W1TO38(-97), .W1TO39(-127), .W1TO40(-111), .W1TO41(-12), .W1TO42(-173), .W1TO43(-13), .W1TO44(-136), .W1TO45(-154), .W1TO46(-81), .W1TO47(-116), .W1TO48(63), .W1TO49(117), .W1TO50(-100), .W1TO51(-80), .W1TO52(-127), .W1TO53(161), .W1TO54(-101), .W1TO55(126), .W1TO56(70), .W1TO57(181), .W1TO58(-145), .W1TO59(22), .W1TO60(76), .W1TO61(137), .W1TO62(143), .W1TO63(105), .W1TO64(58), .W1TO65(41), .W1TO66(73), .W1TO67(-118), .W1TO68(-124), .W1TO69(0), .W1TO70(185), .W1TO71(-28), .W1TO72(100), .W1TO73(-83), .W1TO74(-184), .W1TO75(181), .W1TO76(69), .W1TO77(44), .W1TO78(157), .W1TO79(133), .W1TO80(-143), .W1TO81(-155), .W1TO82(0), .W1TO83(189), .W1TO84(26), .W1TO85(25), .W1TO86(156), .W1TO87(-51), .W1TO88(-100), .W1TO89(186), .W1TO90(133), .W1TO91(-5), .W1TO92(-104), .W1TO93(-80), .W1TO94(148), .W1TO95(74), .W1TO96(-179), .W1TO97(-38), .W1TO98(-13), .W1TO99(-112), .W2TO0(110), .W2TO1(79), .W2TO2(-62), .W2TO3(-77), .W2TO4(89), .W2TO5(126), .W2TO6(171), .W2TO7(8), .W2TO8(-126), .W2TO9(124), .W2TO10(-165), .W2TO11(132), .W2TO12(204), .W2TO13(180), .W2TO14(174), .W2TO15(-153), .W2TO16(-84), .W2TO17(-129), .W2TO18(-116), .W2TO19(-40), .W2TO20(104), .W2TO21(73), .W2TO22(-97), .W2TO23(-39), .W2TO24(-3), .W2TO25(-163), .W2TO26(2), .W2TO27(123), .W2TO28(0), .W2TO29(-14), .W2TO30(-188), .W2TO31(0), .W2TO32(-32), .W2TO33(101), .W2TO34(-176), .W2TO35(125), .W2TO36(15), .W2TO37(4), .W2TO38(127), .W2TO39(36), .W2TO40(-128), .W2TO41(110), .W2TO42(82), .W2TO43(-20), .W2TO44(-27), .W2TO45(90), .W2TO46(139), .W2TO47(-157), .W2TO48(29), .W2TO49(-34), .W2TO50(-80), .W2TO51(-6), .W2TO52(183), .W2TO53(168), .W2TO54(47), .W2TO55(13), .W2TO56(11), .W2TO57(-139), .W2TO58(131), .W2TO59(-74), .W2TO60(-99), .W2TO61(-43), .W2TO62(-51), .W2TO63(137), .W2TO64(58), .W2TO65(3), .W2TO66(141), .W2TO67(-20), .W2TO68(125), .W2TO69(28), .W2TO70(-177), .W2TO71(105), .W2TO72(-168), .W2TO73(49), .W2TO74(-87), .W2TO75(-96), .W2TO76(28), .W2TO77(-94), .W2TO78(-47), .W2TO79(-145), .W2TO80(43), .W2TO81(29), .W2TO82(0), .W2TO83(-26), .W2TO84(-78), .W2TO85(61), .W2TO86(139), .W2TO87(5), .W2TO88(-245), .W2TO89(-67), .W2TO90(14), .W2TO91(-84), .W2TO92(-97), .W2TO93(-77), .W2TO94(77), .W2TO95(38), .W2TO96(194), .W2TO97(145), .W2TO98(-163), .W2TO99(-95), .W3TO0(-99), .W3TO1(-177), .W3TO2(-171), .W3TO3(-57), .W3TO4(170), .W3TO5(-165), .W3TO6(112), .W3TO7(179), .W3TO8(-85), .W3TO9(121), .W3TO10(-88), .W3TO11(-94), .W3TO12(-81), .W3TO13(95), .W3TO14(-171), .W3TO15(-144), .W3TO16(-123), .W3TO17(97), .W3TO18(11), .W3TO19(-181), .W3TO20(-96), .W3TO21(-115), .W3TO22(-147), .W3TO23(-212), .W3TO24(-112), .W3TO25(-91), .W3TO26(-121), .W3TO27(-32), .W3TO28(-37), .W3TO29(2), .W3TO30(-149), .W3TO31(-76), .W3TO32(156), .W3TO33(-93), .W3TO34(72), .W3TO35(105), .W3TO36(121), .W3TO37(-20), .W3TO38(37), .W3TO39(-206), .W3TO40(-220), .W3TO41(-198), .W3TO42(-165), .W3TO43(0), .W3TO44(-127), .W3TO45(-112), .W3TO46(-60), .W3TO47(11), .W3TO48(-17), .W3TO49(44), .W3TO50(173), .W3TO51(-110), .W3TO52(-137), .W3TO53(128), .W3TO54(-48), .W3TO55(-200), .W3TO56(-10), .W3TO57(58), .W3TO58(60), .W3TO59(153), .W3TO60(-215), .W3TO61(29), .W3TO62(-8), .W3TO63(216), .W3TO64(-90), .W3TO65(-144), .W3TO66(53), .W3TO67(-80), .W3TO68(91), .W3TO69(13), .W3TO70(-106), .W3TO71(151), .W3TO72(-3), .W3TO73(-7), .W3TO74(-127), .W3TO75(143), .W3TO76(132), .W3TO77(-46), .W3TO78(49), .W3TO79(154), .W3TO80(-198), .W3TO81(168), .W3TO82(-102), .W3TO83(116), .W3TO84(132), .W3TO85(181), .W3TO86(122), .W3TO87(-196), .W3TO88(-41), .W3TO89(197), .W3TO90(118), .W3TO91(-138), .W3TO92(-143), .W3TO93(-107), .W3TO94(-29), .W3TO95(12), .W3TO96(138), .W3TO97(46), .W3TO98(128), .W3TO99(92), .W4TO0(137), .W4TO1(197), .W4TO2(66), .W4TO3(151), .W4TO4(-40), .W4TO5(16), .W4TO6(202), .W4TO7(-31), .W4TO8(86), .W4TO9(-86), .W4TO10(-65), .W4TO11(59), .W4TO12(46), .W4TO13(-53), .W4TO14(171), .W4TO15(-106), .W4TO16(-148), .W4TO17(-40), .W4TO18(127), .W4TO19(-37), .W4TO20(-142), .W4TO21(-154), .W4TO22(103), .W4TO23(-4), .W4TO24(70), .W4TO25(108), .W4TO26(17), .W4TO27(61), .W4TO28(158), .W4TO29(11), .W4TO30(50), .W4TO31(-122), .W4TO32(-64), .W4TO33(-8), .W4TO34(-15), .W4TO35(42), .W4TO36(-195), .W4TO37(-10), .W4TO38(200), .W4TO39(53), .W4TO40(-241), .W4TO41(90), .W4TO42(-44), .W4TO43(-8), .W4TO44(183), .W4TO45(-174), .W4TO46(-113), .W4TO47(-66), .W4TO48(-110), .W4TO49(126), .W4TO50(2), .W4TO51(12), .W4TO52(0), .W4TO53(181), .W4TO54(-1), .W4TO55(-92), .W4TO56(-58), .W4TO57(-15), .W4TO58(-145), .W4TO59(-12), .W4TO60(-94), .W4TO61(28), .W4TO62(30), .W4TO63(-123), .W4TO64(-30), .W4TO65(143), .W4TO66(5), .W4TO67(-77), .W4TO68(155), .W4TO69(95), .W4TO70(-7), .W4TO71(93), .W4TO72(-41), .W4TO73(-30), .W4TO74(58), .W4TO75(-190), .W4TO76(107), .W4TO77(-60), .W4TO78(-39), .W4TO79(-92), .W4TO80(3), .W4TO81(188), .W4TO82(-105), .W4TO83(159), .W4TO84(-245), .W4TO85(186), .W4TO86(-42), .W4TO87(166), .W4TO88(-131), .W4TO89(-188), .W4TO90(42), .W4TO91(-32), .W4TO92(174), .W4TO93(148), .W4TO94(84), .W4TO95(-111), .W4TO96(148), .W4TO97(-84), .W4TO98(-223), .W4TO99(-12), .W5TO0(-72), .W5TO1(-19), .W5TO2(13), .W5TO3(-30), .W5TO4(-236), .W5TO5(-3), .W5TO6(84), .W5TO7(121), .W5TO8(-48), .W5TO9(137), .W5TO10(158), .W5TO11(106), .W5TO12(86), .W5TO13(1), .W5TO14(41), .W5TO15(-19), .W5TO16(173), .W5TO17(-60), .W5TO18(62), .W5TO19(19), .W5TO20(33), .W5TO21(3), .W5TO22(-46), .W5TO23(-80), .W5TO24(0), .W5TO25(-102), .W5TO26(-124), .W5TO27(-5), .W5TO28(-177), .W5TO29(-290), .W5TO30(-191), .W5TO31(-79), .W5TO32(-113), .W5TO33(32), .W5TO34(-110), .W5TO35(85), .W5TO36(-173), .W5TO37(36), .W5TO38(-21), .W5TO39(-101), .W5TO40(103), .W5TO41(-179), .W5TO42(26), .W5TO43(-51), .W5TO44(-115), .W5TO45(-58), .W5TO46(-5), .W5TO47(120), .W5TO48(63), .W5TO49(-42), .W5TO50(-155), .W5TO51(139), .W5TO52(101), .W5TO53(138), .W5TO54(-35), .W5TO55(138), .W5TO56(-56), .W5TO57(9), .W5TO58(58), .W5TO59(-55), .W5TO60(14), .W5TO61(228), .W5TO62(97), .W5TO63(-34), .W5TO64(8), .W5TO65(138), .W5TO66(-148), .W5TO67(143), .W5TO68(119), .W5TO69(81), .W5TO70(-156), .W5TO71(-30), .W5TO72(99), .W5TO73(-144), .W5TO74(2), .W5TO75(-71), .W5TO76(60), .W5TO77(131), .W5TO78(-36), .W5TO79(236), .W5TO80(66), .W5TO81(-56), .W5TO82(118), .W5TO83(21), .W5TO84(-141), .W5TO85(-100), .W5TO86(-69), .W5TO87(-148), .W5TO88(-65), .W5TO89(196), .W5TO90(182), .W5TO91(-74), .W5TO92(-142), .W5TO93(-143), .W5TO94(-130), .W5TO95(53), .W5TO96(169), .W5TO97(-131), .W5TO98(-36), .W5TO99(157), .W6TO0(19), .W6TO1(-56), .W6TO2(-176), .W6TO3(-98), .W6TO4(-14), .W6TO5(55), .W6TO6(113), .W6TO7(113), .W6TO8(-57), .W6TO9(-162), .W6TO10(-123), .W6TO11(-66), .W6TO12(95), .W6TO13(-75), .W6TO14(-36), .W6TO15(29), .W6TO16(-19), .W6TO17(19), .W6TO18(-66), .W6TO19(-162), .W6TO20(-145), .W6TO21(67), .W6TO22(-23), .W6TO23(-122), .W6TO24(142), .W6TO25(52), .W6TO26(-78), .W6TO27(-33), .W6TO28(-68), .W6TO29(132), .W6TO30(-167), .W6TO31(-184), .W6TO32(0), .W6TO33(-4), .W6TO34(35), .W6TO35(-30), .W6TO36(162), .W6TO37(-1), .W6TO38(61), .W6TO39(-62), .W6TO40(20), .W6TO41(81), .W6TO42(-183), .W6TO43(-67), .W6TO44(60), .W6TO45(60), .W6TO46(7), .W6TO47(89), .W6TO48(-80), .W6TO49(-107), .W6TO50(-106), .W6TO51(145), .W6TO52(55), .W6TO53(-32), .W6TO54(-155), .W6TO55(-189), .W6TO56(-165), .W6TO57(-113), .W6TO58(-183), .W6TO59(29), .W6TO60(-135), .W6TO61(-174), .W6TO62(-86), .W6TO63(-40), .W6TO64(183), .W6TO65(76), .W6TO66(60), .W6TO67(-111), .W6TO68(137), .W6TO69(-72), .W6TO70(-93), .W6TO71(-52), .W6TO72(119), .W6TO73(105), .W6TO74(-188), .W6TO75(141), .W6TO76(-111), .W6TO77(137), .W6TO78(180), .W6TO79(-44), .W6TO80(-207), .W6TO81(1), .W6TO82(-19), .W6TO83(182), .W6TO84(8), .W6TO85(107), .W6TO86(111), .W6TO87(143), .W6TO88(106), .W6TO89(-118), .W6TO90(-125), .W6TO91(12), .W6TO92(93), .W6TO93(68), .W6TO94(-72), .W6TO95(44), .W6TO96(183), .W6TO97(87), .W6TO98(-191), .W6TO99(171), .W7TO0(59), .W7TO1(-151), .W7TO2(-171), .W7TO3(82), .W7TO4(111), .W7TO5(-72), .W7TO6(-47), .W7TO7(99), .W7TO8(-9), .W7TO9(-76), .W7TO10(-58), .W7TO11(-65), .W7TO12(106), .W7TO13(141), .W7TO14(-31), .W7TO15(-133), .W7TO16(79), .W7TO17(-152), .W7TO18(80), .W7TO19(131), .W7TO20(-126), .W7TO21(-119), .W7TO22(-156), .W7TO23(-179), .W7TO24(-84), .W7TO25(91), .W7TO26(-41), .W7TO27(-146), .W7TO28(108), .W7TO29(54), .W7TO30(-151), .W7TO31(177), .W7TO32(137), .W7TO33(-26), .W7TO34(-99), .W7TO35(-65), .W7TO36(88), .W7TO37(139), .W7TO38(-23), .W7TO39(-18), .W7TO40(19), .W7TO41(23), .W7TO42(16), .W7TO43(-12), .W7TO44(126), .W7TO45(30), .W7TO46(55), .W7TO47(105), .W7TO48(36), .W7TO49(-64), .W7TO50(34), .W7TO51(20), .W7TO52(121), .W7TO53(-134), .W7TO54(-187), .W7TO55(-155), .W7TO56(-35), .W7TO57(-82), .W7TO58(46), .W7TO59(65), .W7TO60(36), .W7TO61(157), .W7TO62(-133), .W7TO63(156), .W7TO64(-75), .W7TO65(-47), .W7TO66(-22), .W7TO67(0), .W7TO68(72), .W7TO69(19), .W7TO70(-138), .W7TO71(187), .W7TO72(-13), .W7TO73(29), .W7TO74(130), .W7TO75(16), .W7TO76(-192), .W7TO77(-129), .W7TO78(-1), .W7TO79(-130), .W7TO80(53), .W7TO81(-159), .W7TO82(-134), .W7TO83(8), .W7TO84(146), .W7TO85(-181), .W7TO86(-61), .W7TO87(-62), .W7TO88(-101), .W7TO89(192), .W7TO90(32), .W7TO91(78), .W7TO92(178), .W7TO93(49), .W7TO94(171), .W7TO95(-117), .W7TO96(112), .W7TO97(-46), .W7TO98(-106), .W7TO99(-135), .W8TO0(88), .W8TO1(-159), .W8TO2(26), .W8TO3(124), .W8TO4(-148), .W8TO5(-151), .W8TO6(-91), .W8TO7(-98), .W8TO8(-26), .W8TO9(94), .W8TO10(-188), .W8TO11(-100), .W8TO12(-168), .W8TO13(-82), .W8TO14(159), .W8TO15(114), .W8TO16(-69), .W8TO17(3), .W8TO18(-176), .W8TO19(127), .W8TO20(-64), .W8TO21(-173), .W8TO22(63), .W8TO23(123), .W8TO24(-95), .W8TO25(102), .W8TO26(80), .W8TO27(-6), .W8TO28(-93), .W8TO29(54), .W8TO30(166), .W8TO31(55), .W8TO32(-132), .W8TO33(-107), .W8TO34(67), .W8TO35(45), .W8TO36(73), .W8TO37(25), .W8TO38(76), .W8TO39(-140), .W8TO40(118), .W8TO41(-27), .W8TO42(-170), .W8TO43(-31), .W8TO44(151), .W8TO45(-118), .W8TO46(49), .W8TO47(174), .W8TO48(91), .W8TO49(-155), .W8TO50(-58), .W8TO51(-117), .W8TO52(-54), .W8TO53(184), .W8TO54(-177), .W8TO55(-36), .W8TO56(27), .W8TO57(-118), .W8TO58(175), .W8TO59(127), .W8TO60(80), .W8TO61(174), .W8TO62(-116), .W8TO63(-167), .W8TO64(-86), .W8TO65(127), .W8TO66(20), .W8TO67(-55), .W8TO68(-169), .W8TO69(-10), .W8TO70(109), .W8TO71(111), .W8TO72(-97), .W8TO73(-15), .W8TO74(-73), .W8TO75(-25), .W8TO76(116), .W8TO77(-44), .W8TO78(16), .W8TO79(-32), .W8TO80(-118), .W8TO81(109), .W8TO82(-125), .W8TO83(-57), .W8TO84(111), .W8TO85(131), .W8TO86(-167), .W8TO87(-4), .W8TO88(-105), .W8TO89(-96), .W8TO90(125), .W8TO91(65), .W8TO92(-106), .W8TO93(-58), .W8TO94(184), .W8TO95(34), .W8TO96(175), .W8TO97(-188), .W8TO98(11), .W8TO99(185), .W9TO0(-146), .W9TO1(92), .W9TO2(44), .W9TO3(-108), .W9TO4(-31), .W9TO5(-141), .W9TO6(125), .W9TO7(64), .W9TO8(136), .W9TO9(27), .W9TO10(9), .W9TO11(33), .W9TO12(-58), .W9TO13(-39), .W9TO14(-133), .W9TO15(93), .W9TO16(-71), .W9TO17(-50), .W9TO18(-26), .W9TO19(-107), .W9TO20(-124), .W9TO21(8), .W9TO22(-113), .W9TO23(-119), .W9TO24(74), .W9TO25(-131), .W9TO26(81), .W9TO27(-1), .W9TO28(166), .W9TO29(-138), .W9TO30(-119), .W9TO31(23), .W9TO32(-2), .W9TO33(-72), .W9TO34(90), .W9TO35(-33), .W9TO36(53), .W9TO37(-64), .W9TO38(22), .W9TO39(-191), .W9TO40(-116), .W9TO41(-50), .W9TO42(-37), .W9TO43(84), .W9TO44(-190), .W9TO45(-110), .W9TO46(148), .W9TO47(-71), .W9TO48(-105), .W9TO49(-169), .W9TO50(36), .W9TO51(160), .W9TO52(172), .W9TO53(115), .W9TO54(-74), .W9TO55(-7), .W9TO56(-124), .W9TO57(189), .W9TO58(48), .W9TO59(32), .W9TO60(-133), .W9TO61(-94), .W9TO62(-133), .W9TO63(-48), .W9TO64(112), .W9TO65(-31), .W9TO66(-22), .W9TO67(104), .W9TO68(154), .W9TO69(-24), .W9TO70(-73), .W9TO71(80), .W9TO72(115), .W9TO73(-14), .W9TO74(-131), .W9TO75(-92), .W9TO76(-78), .W9TO77(-113), .W9TO78(-109), .W9TO79(121), .W9TO80(114), .W9TO81(31), .W9TO82(180), .W9TO83(181), .W9TO84(-151), .W9TO85(-171), .W9TO86(5), .W9TO87(-165), .W9TO88(10), .W9TO89(163), .W9TO90(42), .W9TO91(139), .W9TO92(-56), .W9TO93(-140), .W9TO94(-181), .W9TO95(-76), .W9TO96(73), .W9TO97(-159), .W9TO98(-38), .W9TO99(93), .W10TO0(-183), .W10TO1(78), .W10TO2(22), .W10TO3(-168), .W10TO4(4), .W10TO5(73), .W10TO6(-168), .W10TO7(18), .W10TO8(-10), .W10TO9(171), .W10TO10(-199), .W10TO11(-10), .W10TO12(183), .W10TO13(-42), .W10TO14(123), .W10TO15(74), .W10TO16(-123), .W10TO17(31), .W10TO18(153), .W10TO19(-65), .W10TO20(33), .W10TO21(-137), .W10TO22(-4), .W10TO23(34), .W10TO24(258), .W10TO25(-155), .W10TO26(-149), .W10TO27(-27), .W10TO28(29), .W10TO29(69), .W10TO30(94), .W10TO31(0), .W10TO32(-120), .W10TO33(107), .W10TO34(-2), .W10TO35(-53), .W10TO36(77), .W10TO37(14), .W10TO38(-24), .W10TO39(-60), .W10TO40(-7), .W10TO41(-168), .W10TO42(-51), .W10TO43(-30), .W10TO44(23), .W10TO45(133), .W10TO46(-187), .W10TO47(28), .W10TO48(65), .W10TO49(-107), .W10TO50(-42), .W10TO51(29), .W10TO52(63), .W10TO53(-30), .W10TO54(20), .W10TO55(58), .W10TO56(26), .W10TO57(52), .W10TO58(78), .W10TO59(-46), .W10TO60(-251), .W10TO61(-65), .W10TO62(-109), .W10TO63(151), .W10TO64(176), .W10TO65(-159), .W10TO66(-15), .W10TO67(71), .W10TO68(-51), .W10TO69(53), .W10TO70(132), .W10TO71(-137), .W10TO72(94), .W10TO73(-106), .W10TO74(-88), .W10TO75(-189), .W10TO76(20), .W10TO77(-159), .W10TO78(-50), .W10TO79(-91), .W10TO80(75), .W10TO81(-125), .W10TO82(142), .W10TO83(92), .W10TO84(-116), .W10TO85(127), .W10TO86(94), .W10TO87(6), .W10TO88(-126), .W10TO89(-89), .W10TO90(-109), .W10TO91(46), .W10TO92(-29), .W10TO93(-64), .W10TO94(74), .W10TO95(59), .W10TO96(181), .W10TO97(123), .W10TO98(-166), .W10TO99(-37), .W11TO0(-2), .W11TO1(-96), .W11TO2(111), .W11TO3(47), .W11TO4(147), .W11TO5(80), .W11TO6(28), .W11TO7(100), .W11TO8(-112), .W11TO9(21), .W11TO10(143), .W11TO11(135), .W11TO12(141), .W11TO13(-11), .W11TO14(131), .W11TO15(-47), .W11TO16(89), .W11TO17(-62), .W11TO18(-109), .W11TO19(-83), .W11TO20(-144), .W11TO21(58), .W11TO22(-137), .W11TO23(82), .W11TO24(-46), .W11TO25(-115), .W11TO26(-184), .W11TO27(-157), .W11TO28(35), .W11TO29(-19), .W11TO30(181), .W11TO31(83), .W11TO32(44), .W11TO33(126), .W11TO34(-151), .W11TO35(59), .W11TO36(-78), .W11TO37(-4), .W11TO38(187), .W11TO39(68), .W11TO40(-26), .W11TO41(69), .W11TO42(60), .W11TO43(61), .W11TO44(153), .W11TO45(-224), .W11TO46(-113), .W11TO47(51), .W11TO48(-140), .W11TO49(50), .W11TO50(138), .W11TO51(-24), .W11TO52(96), .W11TO53(-61), .W11TO54(5), .W11TO55(160), .W11TO56(-43), .W11TO57(-65), .W11TO58(57), .W11TO59(85), .W11TO60(158), .W11TO61(-104), .W11TO62(-147), .W11TO63(-109), .W11TO64(175), .W11TO65(-85), .W11TO66(-182), .W11TO67(104), .W11TO68(11), .W11TO69(211), .W11TO70(19), .W11TO71(123), .W11TO72(81), .W11TO73(-103), .W11TO74(-83), .W11TO75(21), .W11TO76(-12), .W11TO77(87), .W11TO78(9), .W11TO79(1), .W11TO80(-49), .W11TO81(151), .W11TO82(-109), .W11TO83(10), .W11TO84(53), .W11TO85(16), .W11TO86(-150), .W11TO87(124), .W11TO88(-164), .W11TO89(-81), .W11TO90(-13), .W11TO91(-109), .W11TO92(-1), .W11TO93(3), .W11TO94(-214), .W11TO95(-4), .W11TO96(-45), .W11TO97(-52), .W11TO98(69), .W11TO99(118), .W12TO0(-112), .W12TO1(-67), .W12TO2(61), .W12TO3(42), .W12TO4(38), .W12TO5(-160), .W12TO6(-176), .W12TO7(215), .W12TO8(175), .W12TO9(116), .W12TO10(137), .W12TO11(-92), .W12TO12(150), .W12TO13(45), .W12TO14(-13), .W12TO15(-24), .W12TO16(7), .W12TO17(-38), .W12TO18(-37), .W12TO19(82), .W12TO20(143), .W12TO21(192), .W12TO22(-33), .W12TO23(58), .W12TO24(-63), .W12TO25(-72), .W12TO26(68), .W12TO27(-62), .W12TO28(-155), .W12TO29(18), .W12TO30(-214), .W12TO31(-197), .W12TO32(35), .W12TO33(-158), .W12TO34(72), .W12TO35(-162), .W12TO36(-80), .W12TO37(132), .W12TO38(4), .W12TO39(49), .W12TO40(-139), .W12TO41(-128), .W12TO42(-75), .W12TO43(-184), .W12TO44(113), .W12TO45(-99), .W12TO46(50), .W12TO47(135), .W12TO48(-214), .W12TO49(-40), .W12TO50(47), .W12TO51(5), .W12TO52(151), .W12TO53(24), .W12TO54(-65), .W12TO55(63), .W12TO56(134), .W12TO57(58), .W12TO58(29), .W12TO59(169), .W12TO60(9), .W12TO61(164), .W12TO62(-78), .W12TO63(-131), .W12TO64(-67), .W12TO65(91), .W12TO66(1), .W12TO67(5), .W12TO68(199), .W12TO69(191), .W12TO70(-181), .W12TO71(-109), .W12TO72(-90), .W12TO73(-215), .W12TO74(-126), .W12TO75(174), .W12TO76(31), .W12TO77(-169), .W12TO78(27), .W12TO79(185), .W12TO80(12), .W12TO81(160), .W12TO82(-202), .W12TO83(-18), .W12TO84(-170), .W12TO85(-63), .W12TO86(22), .W12TO87(-45), .W12TO88(-48), .W12TO89(167), .W12TO90(29), .W12TO91(24), .W12TO92(190), .W12TO93(-139), .W12TO94(-198), .W12TO95(-213), .W12TO96(177), .W12TO97(31), .W12TO98(22), .W12TO99(-78), .W13TO0(103), .W13TO1(106), .W13TO2(144), .W13TO3(136), .W13TO4(-52), .W13TO5(90), .W13TO6(-123), .W13TO7(-106), .W13TO8(47), .W13TO9(123), .W13TO10(52), .W13TO11(148), .W13TO12(74), .W13TO13(120), .W13TO14(10), .W13TO15(72), .W13TO16(134), .W13TO17(194), .W13TO18(-202), .W13TO19(73), .W13TO20(-16), .W13TO21(18), .W13TO22(46), .W13TO23(-102), .W13TO24(208), .W13TO25(-138), .W13TO26(94), .W13TO27(123), .W13TO28(-135), .W13TO29(42), .W13TO30(-112), .W13TO31(91), .W13TO32(-30), .W13TO33(141), .W13TO34(-37), .W13TO35(53), .W13TO36(110), .W13TO37(193), .W13TO38(24), .W13TO39(-7), .W13TO40(-54), .W13TO41(0), .W13TO42(-161), .W13TO43(183), .W13TO44(18), .W13TO45(-53), .W13TO46(185), .W13TO47(-27), .W13TO48(-137), .W13TO49(62), .W13TO50(118), .W13TO51(-90), .W13TO52(-105), .W13TO53(-17), .W13TO54(65), .W13TO55(-27), .W13TO56(19), .W13TO57(-180), .W13TO58(-132), .W13TO59(64), .W13TO60(-53), .W13TO61(264), .W13TO62(-136), .W13TO63(-17), .W13TO64(-131), .W13TO65(-187), .W13TO66(96), .W13TO67(-113), .W13TO68(103), .W13TO69(-60), .W13TO70(-82), .W13TO71(-34), .W13TO72(212), .W13TO73(-35), .W13TO74(-176), .W13TO75(-53), .W13TO76(-52), .W13TO77(59), .W13TO78(-8), .W13TO79(233), .W13TO80(49), .W13TO81(-88), .W13TO82(-42), .W13TO83(53), .W13TO84(94), .W13TO85(189), .W13TO86(-168), .W13TO87(75), .W13TO88(68), .W13TO89(153), .W13TO90(-2), .W13TO91(34), .W13TO92(109), .W13TO93(-82), .W13TO94(-146), .W13TO95(-97), .W13TO96(89), .W13TO97(-175), .W13TO98(-107), .W13TO99(88), .W14TO0(-176), .W14TO1(47), .W14TO2(29), .W14TO3(-138), .W14TO4(51), .W14TO5(30), .W14TO6(138), .W14TO7(119), .W14TO8(41), .W14TO9(187), .W14TO10(0), .W14TO11(-64), .W14TO12(61), .W14TO13(116), .W14TO14(71), .W14TO15(-62), .W14TO16(110), .W14TO17(178), .W14TO18(-142), .W14TO19(113), .W14TO20(-146), .W14TO21(94), .W14TO22(-118), .W14TO23(150), .W14TO24(154), .W14TO25(-75), .W14TO26(108), .W14TO27(-178), .W14TO28(-101), .W14TO29(-78), .W14TO30(-71), .W14TO31(-9), .W14TO32(-32), .W14TO33(34), .W14TO34(-74), .W14TO35(25), .W14TO36(-171), .W14TO37(43), .W14TO38(-14), .W14TO39(-86), .W14TO40(-183), .W14TO41(-110), .W14TO42(-26), .W14TO43(11), .W14TO44(-8), .W14TO45(-78), .W14TO46(109), .W14TO47(7), .W14TO48(-7), .W14TO49(46), .W14TO50(-107), .W14TO51(57), .W14TO52(151), .W14TO53(-120), .W14TO54(-40), .W14TO55(118), .W14TO56(190), .W14TO57(123), .W14TO58(114), .W14TO59(73), .W14TO60(-8), .W14TO61(20), .W14TO62(-15), .W14TO63(138), .W14TO64(41), .W14TO65(17), .W14TO66(-175), .W14TO67(63), .W14TO68(-132), .W14TO69(187), .W14TO70(-127), .W14TO71(18), .W14TO72(-155), .W14TO73(-114), .W14TO74(-148), .W14TO75(-130), .W14TO76(-25), .W14TO77(-33), .W14TO78(-101), .W14TO79(53), .W14TO80(-3), .W14TO81(-112), .W14TO82(78), .W14TO83(-128), .W14TO84(102), .W14TO85(-58), .W14TO86(-123), .W14TO87(64), .W14TO88(155), .W14TO89(0), .W14TO90(194), .W14TO91(-164), .W14TO92(-128), .W14TO93(39), .W14TO94(41), .W14TO95(-188), .W14TO96(107), .W14TO97(87), .W14TO98(104), .W14TO99(188), .W15TO0(-152), .W15TO1(-6), .W15TO2(-32), .W15TO3(91), .W15TO4(133), .W15TO5(-35), .W15TO6(30), .W15TO7(133), .W15TO8(-182), .W15TO9(159), .W15TO10(-12), .W15TO11(-65), .W15TO12(93), .W15TO13(153), .W15TO14(-95), .W15TO15(-84), .W15TO16(150), .W15TO17(16), .W15TO18(-72), .W15TO19(-109), .W15TO20(-97), .W15TO21(147), .W15TO22(184), .W15TO23(9), .W15TO24(104), .W15TO25(37), .W15TO26(-55), .W15TO27(28), .W15TO28(-144), .W15TO29(59), .W15TO30(30), .W15TO31(-152), .W15TO32(178), .W15TO33(174), .W15TO34(163), .W15TO35(95), .W15TO36(35), .W15TO37(90), .W15TO38(173), .W15TO39(-174), .W15TO40(20), .W15TO41(-13), .W15TO42(107), .W15TO43(-15), .W15TO44(143), .W15TO45(17), .W15TO46(-20), .W15TO47(-155), .W15TO48(-47), .W15TO49(-109), .W15TO50(89), .W15TO51(-147), .W15TO52(130), .W15TO53(-49), .W15TO54(114), .W15TO55(190), .W15TO56(-140), .W15TO57(-21), .W15TO58(167), .W15TO59(-57), .W15TO60(-167), .W15TO61(119), .W15TO62(63), .W15TO63(-85), .W15TO64(-175), .W15TO65(-95), .W15TO66(160), .W15TO67(129), .W15TO68(141), .W15TO69(-5), .W15TO70(142), .W15TO71(147), .W15TO72(92), .W15TO73(-37), .W15TO74(26), .W15TO75(-169), .W15TO76(-12), .W15TO77(-92), .W15TO78(-183), .W15TO79(-82), .W15TO80(-116), .W15TO81(173), .W15TO82(137), .W15TO83(159), .W15TO84(99), .W15TO85(-124), .W15TO86(-30), .W15TO87(80), .W15TO88(-48), .W15TO89(-66), .W15TO90(-150), .W15TO91(-5), .W15TO92(-105), .W15TO93(-150), .W15TO94(-96), .W15TO95(65), .W15TO96(-106), .W15TO97(-132), .W15TO98(-12), .W15TO99(-27), .W16TO0(-15), .W16TO1(-54), .W16TO2(-189), .W16TO3(25), .W16TO4(-35), .W16TO5(74), .W16TO6(167), .W16TO7(-50), .W16TO8(122), .W16TO9(-122), .W16TO10(93), .W16TO11(-161), .W16TO12(43), .W16TO13(-124), .W16TO14(-147), .W16TO15(-38), .W16TO16(-110), .W16TO17(-127), .W16TO18(136), .W16TO19(121), .W16TO20(164), .W16TO21(-138), .W16TO22(182), .W16TO23(171), .W16TO24(139), .W16TO25(-107), .W16TO26(46), .W16TO27(78), .W16TO28(-8), .W16TO29(151), .W16TO30(125), .W16TO31(70), .W16TO32(-72), .W16TO33(-135), .W16TO34(0), .W16TO35(45), .W16TO36(133), .W16TO37(-34), .W16TO38(-176), .W16TO39(59), .W16TO40(-92), .W16TO41(77), .W16TO42(-48), .W16TO43(9), .W16TO44(173), .W16TO45(-60), .W16TO46(179), .W16TO47(-25), .W16TO48(124), .W16TO49(180), .W16TO50(186), .W16TO51(-164), .W16TO52(168), .W16TO53(26), .W16TO54(104), .W16TO55(42), .W16TO56(111), .W16TO57(-136), .W16TO58(145), .W16TO59(-151), .W16TO60(-40), .W16TO61(15), .W16TO62(-83), .W16TO63(-139), .W16TO64(55), .W16TO65(82), .W16TO66(119), .W16TO67(152), .W16TO68(132), .W16TO69(57), .W16TO70(28), .W16TO71(78), .W16TO72(-149), .W16TO73(-9), .W16TO74(-120), .W16TO75(43), .W16TO76(-131), .W16TO77(-167), .W16TO78(165), .W16TO79(74), .W16TO80(-28), .W16TO81(-24), .W16TO82(-44), .W16TO83(-16), .W16TO84(126), .W16TO85(-13), .W16TO86(146), .W16TO87(158), .W16TO88(-174), .W16TO89(20), .W16TO90(4), .W16TO91(-147), .W16TO92(-97), .W16TO93(110), .W16TO94(41), .W16TO95(134), .W16TO96(-13), .W16TO97(116), .W16TO98(-112), .W16TO99(184), .W17TO0(21), .W17TO1(159), .W17TO2(-152), .W17TO3(143), .W17TO4(-19), .W17TO5(-139), .W17TO6(52), .W17TO7(-207), .W17TO8(103), .W17TO9(134), .W17TO10(-91), .W17TO11(-177), .W17TO12(-50), .W17TO13(79), .W17TO14(-102), .W17TO15(-173), .W17TO16(-36), .W17TO17(179), .W17TO18(-31), .W17TO19(-72), .W17TO20(163), .W17TO21(-8), .W17TO22(200), .W17TO23(138), .W17TO24(125), .W17TO25(-6), .W17TO26(-40), .W17TO27(-21), .W17TO28(0), .W17TO29(73), .W17TO30(-23), .W17TO31(-211), .W17TO32(92), .W17TO33(100), .W17TO34(-115), .W17TO35(38), .W17TO36(24), .W17TO37(-118), .W17TO38(-86), .W17TO39(-126), .W17TO40(161), .W17TO41(39), .W17TO42(164), .W17TO43(-10), .W17TO44(100), .W17TO45(133), .W17TO46(42), .W17TO47(31), .W17TO48(147), .W17TO49(5), .W17TO50(-60), .W17TO51(111), .W17TO52(129), .W17TO53(112), .W17TO54(-156), .W17TO55(30), .W17TO56(-120), .W17TO57(160), .W17TO58(-2), .W17TO59(4), .W17TO60(-116), .W17TO61(-118), .W17TO62(117), .W17TO63(-51), .W17TO64(73), .W17TO65(149), .W17TO66(33), .W17TO67(-116), .W17TO68(171), .W17TO69(171), .W17TO70(41), .W17TO71(-158), .W17TO72(149), .W17TO73(-123), .W17TO74(156), .W17TO75(-69), .W17TO76(-89), .W17TO77(110), .W17TO78(13), .W17TO79(44), .W17TO80(-55), .W17TO81(-130), .W17TO82(-110), .W17TO83(-18), .W17TO84(-77), .W17TO85(-130), .W17TO86(-80), .W17TO87(42), .W17TO88(-51), .W17TO89(0), .W17TO90(-114), .W17TO91(37), .W17TO92(67), .W17TO93(30), .W17TO94(0), .W17TO95(75), .W17TO96(-91), .W17TO97(44), .W17TO98(-142), .W17TO99(-123), .W18TO0(-41), .W18TO1(24), .W18TO2(106), .W18TO3(-108), .W18TO4(159), .W18TO5(43), .W18TO6(128), .W18TO7(-31), .W18TO8(13), .W18TO9(-59), .W18TO10(37), .W18TO11(157), .W18TO12(107), .W18TO13(-62), .W18TO14(-182), .W18TO15(-116), .W18TO16(128), .W18TO17(163), .W18TO18(93), .W18TO19(-133), .W18TO20(99), .W18TO21(149), .W18TO22(-84), .W18TO23(-112), .W18TO24(3), .W18TO25(-121), .W18TO26(-9), .W18TO27(-82), .W18TO28(-173), .W18TO29(-109), .W18TO30(200), .W18TO31(-172), .W18TO32(-40), .W18TO33(19), .W18TO34(-112), .W18TO35(172), .W18TO36(82), .W18TO37(132), .W18TO38(51), .W18TO39(39), .W18TO40(-121), .W18TO41(69), .W18TO42(-158), .W18TO43(63), .W18TO44(-121), .W18TO45(74), .W18TO46(24), .W18TO47(-11), .W18TO48(17), .W18TO49(72), .W18TO50(29), .W18TO51(-62), .W18TO52(106), .W18TO53(-169), .W18TO54(167), .W18TO55(67), .W18TO56(117), .W18TO57(-17), .W18TO58(-113), .W18TO59(61), .W18TO60(33), .W18TO61(-31), .W18TO62(37), .W18TO63(110), .W18TO64(-89), .W18TO65(174), .W18TO66(-62), .W18TO67(-216), .W18TO68(-81), .W18TO69(0), .W18TO70(146), .W18TO71(-123), .W18TO72(-77), .W18TO73(-201), .W18TO74(-182), .W18TO75(-40), .W18TO76(-46), .W18TO77(-92), .W18TO78(-179), .W18TO79(-99), .W18TO80(48), .W18TO81(-59), .W18TO82(143), .W18TO83(76), .W18TO84(197), .W18TO85(-98), .W18TO86(67), .W18TO87(135), .W18TO88(-15), .W18TO89(98), .W18TO90(15), .W18TO91(-55), .W18TO92(191), .W18TO93(-192), .W18TO94(6), .W18TO95(-228), .W18TO96(-32), .W18TO97(61), .W18TO98(124), .W18TO99(47), .W19TO0(-143), .W19TO1(-162), .W19TO2(-87), .W19TO3(160), .W19TO4(-85), .W19TO5(71), .W19TO6(-86), .W19TO7(-131), .W19TO8(52), .W19TO9(-48), .W19TO10(-151), .W19TO11(73), .W19TO12(-11), .W19TO13(-99), .W19TO14(-41), .W19TO15(70), .W19TO16(30), .W19TO17(-41), .W19TO18(-13), .W19TO19(-70), .W19TO20(79), .W19TO21(3), .W19TO22(-34), .W19TO23(-44), .W19TO24(-67), .W19TO25(-40), .W19TO26(-230), .W19TO27(-108), .W19TO28(-109), .W19TO29(-53), .W19TO30(-144), .W19TO31(-14), .W19TO32(118), .W19TO33(-72), .W19TO34(-190), .W19TO35(24), .W19TO36(121), .W19TO37(-63), .W19TO38(70), .W19TO39(107), .W19TO40(-84), .W19TO41(-100), .W19TO42(127), .W19TO43(-123), .W19TO44(105), .W19TO45(-156), .W19TO46(137), .W19TO47(15), .W19TO48(107), .W19TO49(112), .W19TO50(51), .W19TO51(-118), .W19TO52(-82), .W19TO53(61), .W19TO54(112), .W19TO55(159), .W19TO56(-31), .W19TO57(33), .W19TO58(-213), .W19TO59(-22), .W19TO60(220), .W19TO61(-57), .W19TO62(-159), .W19TO63(-80), .W19TO64(32), .W19TO65(193), .W19TO66(-30), .W19TO67(-140), .W19TO68(114), .W19TO69(49), .W19TO70(-154), .W19TO71(-50), .W19TO72(76), .W19TO73(-149), .W19TO74(-184), .W19TO75(-111), .W19TO76(58), .W19TO77(-153), .W19TO78(-17), .W19TO79(92), .W19TO80(57), .W19TO81(24), .W19TO82(53), .W19TO83(-168), .W19TO84(159), .W19TO85(108), .W19TO86(202), .W19TO87(-99), .W19TO88(138), .W19TO89(96), .W19TO90(131), .W19TO91(-95), .W19TO92(57), .W19TO93(-45), .W19TO94(79), .W19TO95(-106), .W19TO96(-79), .W19TO97(147), .W19TO98(177), .W19TO99(69), .W20TO0(26), .W20TO1(50), .W20TO2(-80), .W20TO3(68), .W20TO4(-122), .W20TO5(-27), .W20TO6(55), .W20TO7(-160), .W20TO8(-177), .W20TO9(-121), .W20TO10(163), .W20TO11(-87), .W20TO12(-45), .W20TO13(146), .W20TO14(181), .W20TO15(176), .W20TO16(-207), .W20TO17(170), .W20TO18(171), .W20TO19(179), .W20TO20(-242), .W20TO21(-93), .W20TO22(-27), .W20TO23(-121), .W20TO24(-119), .W20TO25(26), .W20TO26(-41), .W20TO27(-142), .W20TO28(-28), .W20TO29(-89), .W20TO30(0), .W20TO31(-50), .W20TO32(32), .W20TO33(27), .W20TO34(135), .W20TO35(-11), .W20TO36(-149), .W20TO37(108), .W20TO38(74), .W20TO39(-75), .W20TO40(-25), .W20TO41(17), .W20TO42(-170), .W20TO43(139), .W20TO44(-150), .W20TO45(-207), .W20TO46(-147), .W20TO47(275), .W20TO48(-188), .W20TO49(-124), .W20TO50(-136), .W20TO51(-101), .W20TO52(-142), .W20TO53(50), .W20TO54(46), .W20TO55(13), .W20TO56(-83), .W20TO57(61), .W20TO58(41), .W20TO59(-205), .W20TO60(73), .W20TO61(-36), .W20TO62(-32), .W20TO63(0), .W20TO64(-137), .W20TO65(53), .W20TO66(-75), .W20TO67(-116), .W20TO68(-114), .W20TO69(19), .W20TO70(26), .W20TO71(-84), .W20TO72(161), .W20TO73(114), .W20TO74(-135), .W20TO75(-89), .W20TO76(106), .W20TO77(189), .W20TO78(114), .W20TO79(-61), .W20TO80(-124), .W20TO81(133), .W20TO82(1), .W20TO83(-75), .W20TO84(27), .W20TO85(-37), .W20TO86(80), .W20TO87(-228), .W20TO88(-44), .W20TO89(62), .W20TO90(130), .W20TO91(144), .W20TO92(3), .W20TO93(16), .W20TO94(-29), .W20TO95(80), .W20TO96(53), .W20TO97(-32), .W20TO98(70), .W20TO99(39), .W21TO0(-119), .W21TO1(49), .W21TO2(65), .W21TO3(-187), .W21TO4(111), .W21TO5(-335), .W21TO6(-38), .W21TO7(-79), .W21TO8(-58), .W21TO9(48), .W21TO10(-94), .W21TO11(200), .W21TO12(42), .W21TO13(141), .W21TO14(-2), .W21TO15(210), .W21TO16(-44), .W21TO17(-103), .W21TO18(-157), .W21TO19(15), .W21TO20(-220), .W21TO21(125), .W21TO22(172), .W21TO23(95), .W21TO24(170), .W21TO25(149), .W21TO26(-183), .W21TO27(-57), .W21TO28(-93), .W21TO29(119), .W21TO30(-17), .W21TO31(-78), .W21TO32(-28), .W21TO33(-251), .W21TO34(99), .W21TO35(18), .W21TO36(-186), .W21TO37(189), .W21TO38(91), .W21TO39(-46), .W21TO40(121), .W21TO41(102), .W21TO42(-93), .W21TO43(-32), .W21TO44(-175), .W21TO45(74), .W21TO46(-99), .W21TO47(245), .W21TO48(-151), .W21TO49(-93), .W21TO50(162), .W21TO51(85), .W21TO52(95), .W21TO53(-253), .W21TO54(-191), .W21TO55(-31), .W21TO56(-131), .W21TO57(-26), .W21TO58(137), .W21TO59(-40), .W21TO60(-5), .W21TO61(130), .W21TO62(-155), .W21TO63(175), .W21TO64(-32), .W21TO65(-79), .W21TO66(101), .W21TO67(-77), .W21TO68(113), .W21TO69(138), .W21TO70(163), .W21TO71(211), .W21TO72(-60), .W21TO73(130), .W21TO74(118), .W21TO75(72), .W21TO76(-173), .W21TO77(-109), .W21TO78(-35), .W21TO79(-172), .W21TO80(147), .W21TO81(2), .W21TO82(9), .W21TO83(-30), .W21TO84(28), .W21TO85(-43), .W21TO86(83), .W21TO87(59), .W21TO88(0), .W21TO89(67), .W21TO90(23), .W21TO91(-30), .W21TO92(-3), .W21TO93(2), .W21TO94(10), .W21TO95(17), .W21TO96(-73), .W21TO97(-129), .W21TO98(110), .W21TO99(136), .W22TO0(-65), .W22TO1(57), .W22TO2(-123), .W22TO3(-192), .W22TO4(-152), .W22TO5(-136), .W22TO6(65), .W22TO7(-104), .W22TO8(-53), .W22TO9(-48), .W22TO10(189), .W22TO11(37), .W22TO12(-154), .W22TO13(113), .W22TO14(186), .W22TO15(-156), .W22TO16(75), .W22TO17(-97), .W22TO18(-185), .W22TO19(-102), .W22TO20(5), .W22TO21(-161), .W22TO22(139), .W22TO23(67), .W22TO24(-62), .W22TO25(-94), .W22TO26(-84), .W22TO27(111), .W22TO28(9), .W22TO29(67), .W22TO30(137), .W22TO31(-102), .W22TO32(204), .W22TO33(101), .W22TO34(57), .W22TO35(32), .W22TO36(0), .W22TO37(115), .W22TO38(-44), .W22TO39(101), .W22TO40(-138), .W22TO41(197), .W22TO42(17), .W22TO43(173), .W22TO44(-33), .W22TO45(-43), .W22TO46(78), .W22TO47(145), .W22TO48(-147), .W22TO49(104), .W22TO50(-65), .W22TO51(-97), .W22TO52(70), .W22TO53(-96), .W22TO54(-54), .W22TO55(81), .W22TO56(-127), .W22TO57(97), .W22TO58(-86), .W22TO59(89), .W22TO60(-37), .W22TO61(220), .W22TO62(-188), .W22TO63(35), .W22TO64(174), .W22TO65(-90), .W22TO66(-35), .W22TO67(-91), .W22TO68(104), .W22TO69(190), .W22TO70(-17), .W22TO71(0), .W22TO72(-101), .W22TO73(126), .W22TO74(-141), .W22TO75(-69), .W22TO76(122), .W22TO77(-179), .W22TO78(39), .W22TO79(-59), .W22TO80(-88), .W22TO81(147), .W22TO82(11), .W22TO83(-136), .W22TO84(136), .W22TO85(-107), .W22TO86(120), .W22TO87(-113), .W22TO88(-28), .W22TO89(105), .W22TO90(71), .W22TO91(23), .W22TO92(88), .W22TO93(-91), .W22TO94(-152), .W22TO95(113), .W22TO96(179), .W22TO97(-176), .W22TO98(-27), .W22TO99(-9), .W23TO0(-157), .W23TO1(101), .W23TO2(155), .W23TO3(-37), .W23TO4(-182), .W23TO5(-13), .W23TO6(88), .W23TO7(-62), .W23TO8(109), .W23TO9(-50), .W23TO10(125), .W23TO11(-57), .W23TO12(-123), .W23TO13(-53), .W23TO14(30), .W23TO15(-151), .W23TO16(-145), .W23TO17(-19), .W23TO18(-71), .W23TO19(-98), .W23TO20(-24), .W23TO21(-2), .W23TO22(24), .W23TO23(152), .W23TO24(-12), .W23TO25(-22), .W23TO26(-101), .W23TO27(72), .W23TO28(-188), .W23TO29(-119), .W23TO30(-44), .W23TO31(151), .W23TO32(118), .W23TO33(-120), .W23TO34(185), .W23TO35(-53), .W23TO36(-34), .W23TO37(185), .W23TO38(143), .W23TO39(-123), .W23TO40(24), .W23TO41(-87), .W23TO42(-140), .W23TO43(-9), .W23TO44(-9), .W23TO45(151), .W23TO46(142), .W23TO47(-169), .W23TO48(9), .W23TO49(26), .W23TO50(-96), .W23TO51(-121), .W23TO52(18), .W23TO53(170), .W23TO54(-39), .W23TO55(-73), .W23TO56(69), .W23TO57(52), .W23TO58(-59), .W23TO59(65), .W23TO60(-119), .W23TO61(47), .W23TO62(-117), .W23TO63(147), .W23TO64(111), .W23TO65(97), .W23TO66(123), .W23TO67(-68), .W23TO68(123), .W23TO69(-82), .W23TO70(30), .W23TO71(93), .W23TO72(-126), .W23TO73(-179), .W23TO74(18), .W23TO75(-103), .W23TO76(154), .W23TO77(177), .W23TO78(-43), .W23TO79(174), .W23TO80(-11), .W23TO81(-91), .W23TO82(-34), .W23TO83(133), .W23TO84(6), .W23TO85(-44), .W23TO86(69), .W23TO87(-73), .W23TO88(-120), .W23TO89(119), .W23TO90(-35), .W23TO91(-56), .W23TO92(185), .W23TO93(189), .W23TO94(73), .W23TO95(122), .W23TO96(67), .W23TO97(-21), .W23TO98(-104), .W23TO99(5), .W24TO0(-185), .W24TO1(5), .W24TO2(47), .W24TO3(10), .W24TO4(-29), .W24TO5(-121), .W24TO6(54), .W24TO7(-48), .W24TO8(105), .W24TO9(-179), .W24TO10(-155), .W24TO11(149), .W24TO12(-94), .W24TO13(-95), .W24TO14(-184), .W24TO15(-27), .W24TO16(15), .W24TO17(16), .W24TO18(186), .W24TO19(-135), .W24TO20(-141), .W24TO21(-30), .W24TO22(30), .W24TO23(20), .W24TO24(99), .W24TO25(-32), .W24TO26(-40), .W24TO27(74), .W24TO28(-188), .W24TO29(72), .W24TO30(82), .W24TO31(169), .W24TO32(74), .W24TO33(-16), .W24TO34(-175), .W24TO35(7), .W24TO36(-177), .W24TO37(163), .W24TO38(102), .W24TO39(-11), .W24TO40(-116), .W24TO41(79), .W24TO42(-31), .W24TO43(-58), .W24TO44(-32), .W24TO45(35), .W24TO46(51), .W24TO47(165), .W24TO48(-140), .W24TO49(-17), .W24TO50(81), .W24TO51(80), .W24TO52(163), .W24TO53(-46), .W24TO54(186), .W24TO55(-112), .W24TO56(56), .W24TO57(168), .W24TO58(53), .W24TO59(94), .W24TO60(-61), .W24TO61(-179), .W24TO62(-106), .W24TO63(-66), .W24TO64(-117), .W24TO65(-63), .W24TO66(114), .W24TO67(-63), .W24TO68(-5), .W24TO69(149), .W24TO70(144), .W24TO71(-114), .W24TO72(99), .W24TO73(-19), .W24TO74(26), .W24TO75(91), .W24TO76(47), .W24TO77(168), .W24TO78(115), .W24TO79(-82), .W24TO80(-14), .W24TO81(-123), .W24TO82(-73), .W24TO83(120), .W24TO84(-100), .W24TO85(-187), .W24TO86(135), .W24TO87(-7), .W24TO88(149), .W24TO89(186), .W24TO90(0), .W24TO91(-43), .W24TO92(-131), .W24TO93(-90), .W24TO94(-149), .W24TO95(-94), .W24TO96(-56), .W24TO97(-191), .W24TO98(6), .W24TO99(153), .W25TO0(-160), .W25TO1(132), .W25TO2(-7), .W25TO3(111), .W25TO4(-202), .W25TO5(116), .W25TO6(86), .W25TO7(23), .W25TO8(-126), .W25TO9(-75), .W25TO10(-22), .W25TO11(94), .W25TO12(141), .W25TO13(-189), .W25TO14(19), .W25TO15(-44), .W25TO16(183), .W25TO17(33), .W25TO18(-32), .W25TO19(-93), .W25TO20(179), .W25TO21(1), .W25TO22(-82), .W25TO23(76), .W25TO24(-121), .W25TO25(-28), .W25TO26(-110), .W25TO27(160), .W25TO28(-159), .W25TO29(-78), .W25TO30(-117), .W25TO31(91), .W25TO32(45), .W25TO33(19), .W25TO34(-8), .W25TO35(-144), .W25TO36(160), .W25TO37(-75), .W25TO38(92), .W25TO39(-31), .W25TO40(83), .W25TO41(68), .W25TO42(-180), .W25TO43(-90), .W25TO44(-108), .W25TO45(-151), .W25TO46(-72), .W25TO47(-120), .W25TO48(-161), .W25TO49(-117), .W25TO50(-189), .W25TO51(126), .W25TO52(-188), .W25TO53(-124), .W25TO54(-48), .W25TO55(-50), .W25TO56(194), .W25TO57(4), .W25TO58(-133), .W25TO59(71), .W25TO60(91), .W25TO61(29), .W25TO62(88), .W25TO63(-89), .W25TO64(-22), .W25TO65(-102), .W25TO66(-178), .W25TO67(-35), .W25TO68(-68), .W25TO69(117), .W25TO70(81), .W25TO71(48), .W25TO72(67), .W25TO73(47), .W25TO74(-52), .W25TO75(0), .W25TO76(193), .W25TO77(-198), .W25TO78(101), .W25TO79(-142), .W25TO80(-8), .W25TO81(-51), .W25TO82(-179), .W25TO83(64), .W25TO84(6), .W25TO85(-90), .W25TO86(127), .W25TO87(147), .W25TO88(-71), .W25TO89(-164), .W25TO90(82), .W25TO91(134), .W25TO92(63), .W25TO93(5), .W25TO94(-81), .W25TO95(-193), .W25TO96(54), .W25TO97(178), .W25TO98(92), .W25TO99(-39), .W26TO0(-124), .W26TO1(-20), .W26TO2(-121), .W26TO3(164), .W26TO4(30), .W26TO5(151), .W26TO6(113), .W26TO7(-237), .W26TO8(-145), .W26TO9(150), .W26TO10(131), .W26TO11(140), .W26TO12(-89), .W26TO13(-25), .W26TO14(158), .W26TO15(26), .W26TO16(157), .W26TO17(-67), .W26TO18(-119), .W26TO19(-197), .W26TO20(-59), .W26TO21(-143), .W26TO22(111), .W26TO23(-153), .W26TO24(-259), .W26TO25(58), .W26TO26(71), .W26TO27(-43), .W26TO28(-107), .W26TO29(128), .W26TO30(-107), .W26TO31(42), .W26TO32(46), .W26TO33(-27), .W26TO34(-46), .W26TO35(64), .W26TO36(-28), .W26TO37(-56), .W26TO38(-153), .W26TO39(93), .W26TO40(-55), .W26TO41(3), .W26TO42(86), .W26TO43(79), .W26TO44(115), .W26TO45(-156), .W26TO46(-41), .W26TO47(-81), .W26TO48(44), .W26TO49(192), .W26TO50(-134), .W26TO51(-36), .W26TO52(86), .W26TO53(-69), .W26TO54(175), .W26TO55(-198), .W26TO56(-38), .W26TO57(28), .W26TO58(36), .W26TO59(-241), .W26TO60(144), .W26TO61(-143), .W26TO62(-123), .W26TO63(67), .W26TO64(-85), .W26TO65(-99), .W26TO66(-207), .W26TO67(-94), .W26TO68(7), .W26TO69(32), .W26TO70(-195), .W26TO71(110), .W26TO72(-70), .W26TO73(61), .W26TO74(62), .W26TO75(43), .W26TO76(-145), .W26TO77(95), .W26TO78(80), .W26TO79(-204), .W26TO80(-36), .W26TO81(171), .W26TO82(61), .W26TO83(-166), .W26TO84(-106), .W26TO85(125), .W26TO86(63), .W26TO87(102), .W26TO88(78), .W26TO89(-127), .W26TO90(188), .W26TO91(-299), .W26TO92(102), .W26TO93(-258), .W26TO94(-106), .W26TO95(-136), .W26TO96(-6), .W26TO97(-33), .W26TO98(34), .W26TO99(-84), .W27TO0(-64), .W27TO1(80), .W27TO2(-47), .W27TO3(-52), .W27TO4(-125), .W27TO5(-86), .W27TO6(96), .W27TO7(12), .W27TO8(226), .W27TO9(-65), .W27TO10(166), .W27TO11(-140), .W27TO12(137), .W27TO13(129), .W27TO14(-190), .W27TO15(12), .W27TO16(-73), .W27TO17(46), .W27TO18(-28), .W27TO19(65), .W27TO20(-83), .W27TO21(139), .W27TO22(69), .W27TO23(-14), .W27TO24(-47), .W27TO25(148), .W27TO26(-27), .W27TO27(42), .W27TO28(-68), .W27TO29(-121), .W27TO30(94), .W27TO31(56), .W27TO32(-113), .W27TO33(-14), .W27TO34(-118), .W27TO35(63), .W27TO36(32), .W27TO37(45), .W27TO38(-177), .W27TO39(64), .W27TO40(-44), .W27TO41(-24), .W27TO42(110), .W27TO43(-43), .W27TO44(99), .W27TO45(-7), .W27TO46(-112), .W27TO47(9), .W27TO48(114), .W27TO49(157), .W27TO50(-91), .W27TO51(24), .W27TO52(-160), .W27TO53(-100), .W27TO54(-129), .W27TO55(152), .W27TO56(9), .W27TO57(-60), .W27TO58(-226), .W27TO59(-273), .W27TO60(-30), .W27TO61(-75), .W27TO62(132), .W27TO63(172), .W27TO64(-72), .W27TO65(-47), .W27TO66(55), .W27TO67(25), .W27TO68(164), .W27TO69(-64), .W27TO70(118), .W27TO71(175), .W27TO72(-129), .W27TO73(34), .W27TO74(165), .W27TO75(-146), .W27TO76(-69), .W27TO77(-135), .W27TO78(-271), .W27TO79(-26), .W27TO80(31), .W27TO81(-32), .W27TO82(166), .W27TO83(22), .W27TO84(222), .W27TO85(108), .W27TO86(28), .W27TO87(176), .W27TO88(182), .W27TO89(-119), .W27TO90(-38), .W27TO91(-47), .W27TO92(-126), .W27TO93(-35), .W27TO94(-3), .W27TO95(-104), .W27TO96(106), .W27TO97(-79), .W27TO98(-154), .W27TO99(-54), .W28TO0(-48), .W28TO1(-58), .W28TO2(-283), .W28TO3(-205), .W28TO4(-211), .W28TO5(36), .W28TO6(-6), .W28TO7(45), .W28TO8(-113), .W28TO9(-3), .W28TO10(-166), .W28TO11(95), .W28TO12(150), .W28TO13(72), .W28TO14(-81), .W28TO15(55), .W28TO16(146), .W28TO17(30), .W28TO18(216), .W28TO19(-144), .W28TO20(131), .W28TO21(-168), .W28TO22(-91), .W28TO23(139), .W28TO24(-129), .W28TO25(96), .W28TO26(-97), .W28TO27(-106), .W28TO28(44), .W28TO29(133), .W28TO30(-43), .W28TO31(-25), .W28TO32(10), .W28TO33(-118), .W28TO34(23), .W28TO35(93), .W28TO36(39), .W28TO37(78), .W28TO38(-129), .W28TO39(-113), .W28TO40(32), .W28TO41(-151), .W28TO42(69), .W28TO43(-149), .W28TO44(79), .W28TO45(46), .W28TO46(-127), .W28TO47(72), .W28TO48(134), .W28TO49(100), .W28TO50(36), .W28TO51(-150), .W28TO52(-80), .W28TO53(165), .W28TO54(-125), .W28TO55(-82), .W28TO56(153), .W28TO57(104), .W28TO58(65), .W28TO59(-65), .W28TO60(-18), .W28TO61(98), .W28TO62(40), .W28TO63(-26), .W28TO64(37), .W28TO65(40), .W28TO66(-48), .W28TO67(-43), .W28TO68(93), .W28TO69(0), .W28TO70(-28), .W28TO71(101), .W28TO72(-102), .W28TO73(-205), .W28TO74(15), .W28TO75(-115), .W28TO76(-87), .W28TO77(-26), .W28TO78(-96), .W28TO79(68), .W28TO80(-165), .W28TO81(160), .W28TO82(252), .W28TO83(36), .W28TO84(1), .W28TO85(-48), .W28TO86(-85), .W28TO87(26), .W28TO88(41), .W28TO89(87), .W28TO90(79), .W28TO91(-40), .W28TO92(161), .W28TO93(54), .W28TO94(-32), .W28TO95(263), .W28TO96(-108), .W28TO97(33), .W28TO98(77), .W28TO99(-60), .W29TO0(-120), .W29TO1(-58), .W29TO2(194), .W29TO3(-54), .W29TO4(-118), .W29TO5(-64), .W29TO6(147), .W29TO7(19), .W29TO8(-59), .W29TO9(53), .W29TO10(132), .W29TO11(-5), .W29TO12(0), .W29TO13(172), .W29TO14(-161), .W29TO15(176), .W29TO16(255), .W29TO17(-58), .W29TO18(-24), .W29TO19(-17), .W29TO20(31), .W29TO21(58), .W29TO22(164), .W29TO23(-133), .W29TO24(-134), .W29TO25(24), .W29TO26(25), .W29TO27(-168), .W29TO28(-27), .W29TO29(173), .W29TO30(-46), .W29TO31(-124), .W29TO32(70), .W29TO33(-1), .W29TO34(-81), .W29TO35(-15), .W29TO36(-136), .W29TO37(40), .W29TO38(94), .W29TO39(88), .W29TO40(16), .W29TO41(-129), .W29TO42(160), .W29TO43(-11), .W29TO44(-40), .W29TO45(-185), .W29TO46(-5), .W29TO47(92), .W29TO48(139), .W29TO49(115), .W29TO50(38), .W29TO51(128), .W29TO52(123), .W29TO53(-123), .W29TO54(4), .W29TO55(-42), .W29TO56(69), .W29TO57(-133), .W29TO58(-39), .W29TO59(-119), .W29TO60(-55), .W29TO61(-96), .W29TO62(-111), .W29TO63(-64), .W29TO64(-132), .W29TO65(153), .W29TO66(70), .W29TO67(-220), .W29TO68(-35), .W29TO69(-74), .W29TO70(-5), .W29TO71(-69), .W29TO72(170), .W29TO73(-25), .W29TO74(31), .W29TO75(-21), .W29TO76(-237), .W29TO77(57), .W29TO78(73), .W29TO79(-126), .W29TO80(33), .W29TO81(-76), .W29TO82(-238), .W29TO83(-29), .W29TO84(209), .W29TO85(209), .W29TO86(-19), .W29TO87(-90), .W29TO88(-101), .W29TO89(-126), .W29TO90(-65), .W29TO91(-133), .W29TO92(201), .W29TO93(-41), .W29TO94(-214), .W29TO95(-203), .W29TO96(-136), .W29TO97(-162), .W29TO98(96), .W29TO99(170), .W30TO0(-25), .W30TO1(-68), .W30TO2(92), .W30TO3(77), .W30TO4(123), .W30TO5(0), .W30TO6(64), .W30TO7(-60), .W30TO8(-32), .W30TO9(182), .W30TO10(-144), .W30TO11(-108), .W30TO12(76), .W30TO13(-100), .W30TO14(191), .W30TO15(-172), .W30TO16(91), .W30TO17(140), .W30TO18(66), .W30TO19(-179), .W30TO20(-174), .W30TO21(-36), .W30TO22(10), .W30TO23(124), .W30TO24(102), .W30TO25(-163), .W30TO26(-59), .W30TO27(48), .W30TO28(-89), .W30TO29(249), .W30TO30(-3), .W30TO31(143), .W30TO32(18), .W30TO33(-95), .W30TO34(47), .W30TO35(28), .W30TO36(14), .W30TO37(-31), .W30TO38(85), .W30TO39(-71), .W30TO40(-182), .W30TO41(21), .W30TO42(20), .W30TO43(-103), .W30TO44(123), .W30TO45(115), .W30TO46(-186), .W30TO47(-144), .W30TO48(164), .W30TO49(101), .W30TO50(133), .W30TO51(163), .W30TO52(-90), .W30TO53(-65), .W30TO54(188), .W30TO55(-34), .W30TO56(-19), .W30TO57(25), .W30TO58(-11), .W30TO59(-184), .W30TO60(44), .W30TO61(32), .W30TO62(156), .W30TO63(-130), .W30TO64(55), .W30TO65(62), .W30TO66(-84), .W30TO67(-112), .W30TO68(118), .W30TO69(39), .W30TO70(99), .W30TO71(115), .W30TO72(56), .W30TO73(-94), .W30TO74(-82), .W30TO75(128), .W30TO76(-7), .W30TO77(145), .W30TO78(212), .W30TO79(-17), .W30TO80(88), .W30TO81(-8), .W30TO82(-220), .W30TO83(86), .W30TO84(63), .W30TO85(165), .W30TO86(135), .W30TO87(137), .W30TO88(-74), .W30TO89(-90), .W30TO90(168), .W30TO91(-52), .W30TO92(190), .W30TO93(-57), .W30TO94(100), .W30TO95(4), .W30TO96(13), .W30TO97(-133), .W30TO98(150), .W30TO99(-180), .W31TO0(-65), .W31TO1(-106), .W31TO2(-155), .W31TO3(59), .W31TO4(141), .W31TO5(-59), .W31TO6(-22), .W31TO7(72), .W31TO8(-70), .W31TO9(-157), .W31TO10(14), .W31TO11(156), .W31TO12(0), .W31TO13(104), .W31TO14(54), .W31TO15(-21), .W31TO16(4), .W31TO17(-155), .W31TO18(-174), .W31TO19(-119), .W31TO20(-178), .W31TO21(-70), .W31TO22(-55), .W31TO23(-149), .W31TO24(56), .W31TO25(80), .W31TO26(-31), .W31TO27(-101), .W31TO28(-15), .W31TO29(-60), .W31TO30(-29), .W31TO31(77), .W31TO32(15), .W31TO33(88), .W31TO34(-163), .W31TO35(88), .W31TO36(106), .W31TO37(146), .W31TO38(149), .W31TO39(53), .W31TO40(-68), .W31TO41(56), .W31TO42(-113), .W31TO43(91), .W31TO44(35), .W31TO45(43), .W31TO46(-123), .W31TO47(-27), .W31TO48(-96), .W31TO49(-83), .W31TO50(184), .W31TO51(0), .W31TO52(-154), .W31TO53(-152), .W31TO54(148), .W31TO55(-125), .W31TO56(3), .W31TO57(40), .W31TO58(-189), .W31TO59(-89), .W31TO60(-137), .W31TO61(-97), .W31TO62(-181), .W31TO63(148), .W31TO64(98), .W31TO65(42), .W31TO66(161), .W31TO67(140), .W31TO68(-40), .W31TO69(102), .W31TO70(125), .W31TO71(176), .W31TO72(37), .W31TO73(-33), .W31TO74(111), .W31TO75(-176), .W31TO76(-96), .W31TO77(28), .W31TO78(-173), .W31TO79(154), .W31TO80(-151), .W31TO81(165), .W31TO82(186), .W31TO83(-117), .W31TO84(-40), .W31TO85(91), .W31TO86(157), .W31TO87(169), .W31TO88(-185), .W31TO89(-107), .W31TO90(87), .W31TO91(3), .W31TO92(113), .W31TO93(-72), .W31TO94(116), .W31TO95(84), .W31TO96(-77), .W31TO97(-187), .W31TO98(-77), .W31TO99(-63), .W32TO0(90), .W32TO1(-112), .W32TO2(-112), .W32TO3(-59), .W32TO4(-145), .W32TO5(127), .W32TO6(-178), .W32TO7(-189), .W32TO8(-64), .W32TO9(-79), .W32TO10(186), .W32TO11(0), .W32TO12(-39), .W32TO13(141), .W32TO14(59), .W32TO15(-2), .W32TO16(-167), .W32TO17(14), .W32TO18(92), .W32TO19(138), .W32TO20(-109), .W32TO21(50), .W32TO22(168), .W32TO23(102), .W32TO24(107), .W32TO25(-4), .W32TO26(-3), .W32TO27(-120), .W32TO28(34), .W32TO29(-65), .W32TO30(27), .W32TO31(-69), .W32TO32(-188), .W32TO33(108), .W32TO34(-61), .W32TO35(-116), .W32TO36(157), .W32TO37(-93), .W32TO38(-176), .W32TO39(162), .W32TO40(-158), .W32TO41(-58), .W32TO42(99), .W32TO43(-140), .W32TO44(-172), .W32TO45(-102), .W32TO46(-41), .W32TO47(-149), .W32TO48(-43), .W32TO49(-50), .W32TO50(154), .W32TO51(-15), .W32TO52(-10), .W32TO53(159), .W32TO54(-151), .W32TO55(-136), .W32TO56(158), .W32TO57(-105), .W32TO58(-172), .W32TO59(-64), .W32TO60(75), .W32TO61(-124), .W32TO62(-177), .W32TO63(77), .W32TO64(-103), .W32TO65(-8), .W32TO66(156), .W32TO67(-111), .W32TO68(-118), .W32TO69(125), .W32TO70(110), .W32TO71(-141), .W32TO72(-186), .W32TO73(95), .W32TO74(-80), .W32TO75(-62), .W32TO76(96), .W32TO77(72), .W32TO78(102), .W32TO79(-129), .W32TO80(-38), .W32TO81(37), .W32TO82(19), .W32TO83(186), .W32TO84(-26), .W32TO85(27), .W32TO86(105), .W32TO87(72), .W32TO88(-121), .W32TO89(35), .W32TO90(-164), .W32TO91(144), .W32TO92(-37), .W32TO93(-102), .W32TO94(100), .W32TO95(179), .W32TO96(-82), .W32TO97(-24), .W32TO98(-138), .W32TO99(11), .W33TO0(174), .W33TO1(-126), .W33TO2(114), .W33TO3(-32), .W33TO4(-49), .W33TO5(-134), .W33TO6(-124), .W33TO7(-130), .W33TO8(104), .W33TO9(58), .W33TO10(171), .W33TO11(-120), .W33TO12(76), .W33TO13(-210), .W33TO14(-145), .W33TO15(59), .W33TO16(-59), .W33TO17(163), .W33TO18(-135), .W33TO19(-120), .W33TO20(-151), .W33TO21(-19), .W33TO22(-222), .W33TO23(6), .W33TO24(-139), .W33TO25(-68), .W33TO26(-84), .W33TO27(-181), .W33TO28(-1), .W33TO29(112), .W33TO30(-132), .W33TO31(-84), .W33TO32(-156), .W33TO33(28), .W33TO34(115), .W33TO35(-63), .W33TO36(-75), .W33TO37(16), .W33TO38(180), .W33TO39(19), .W33TO40(24), .W33TO41(14), .W33TO42(54), .W33TO43(-133), .W33TO44(-183), .W33TO45(-2), .W33TO46(-137), .W33TO47(-196), .W33TO48(111), .W33TO49(135), .W33TO50(26), .W33TO51(-139), .W33TO52(17), .W33TO53(-104), .W33TO54(54), .W33TO55(30), .W33TO56(177), .W33TO57(76), .W33TO58(-92), .W33TO59(124), .W33TO60(86), .W33TO61(95), .W33TO62(-60), .W33TO63(-184), .W33TO64(-64), .W33TO65(-63), .W33TO66(-133), .W33TO67(-118), .W33TO68(-83), .W33TO69(100), .W33TO70(-204), .W33TO71(-74), .W33TO72(-99), .W33TO73(-110), .W33TO74(-3), .W33TO75(173), .W33TO76(79), .W33TO77(-162), .W33TO78(6), .W33TO79(-164), .W33TO80(-71), .W33TO81(-49), .W33TO82(-273), .W33TO83(-199), .W33TO84(-6), .W33TO85(99), .W33TO86(-58), .W33TO87(172), .W33TO88(-41), .W33TO89(93), .W33TO90(-173), .W33TO91(103), .W33TO92(-96), .W33TO93(64), .W33TO94(-200), .W33TO95(-89), .W33TO96(25), .W33TO97(-143), .W33TO98(-31), .W33TO99(-180), .W34TO0(-60), .W34TO1(-30), .W34TO2(-163), .W34TO3(-182), .W34TO4(92), .W34TO5(-105), .W34TO6(-157), .W34TO7(-9), .W34TO8(216), .W34TO9(116), .W34TO10(95), .W34TO11(14), .W34TO12(27), .W34TO13(-108), .W34TO14(-183), .W34TO15(-11), .W34TO16(94), .W34TO17(-153), .W34TO18(33), .W34TO19(-124), .W34TO20(-50), .W34TO21(-143), .W34TO22(-226), .W34TO23(80), .W34TO24(-222), .W34TO25(-210), .W34TO26(132), .W34TO27(37), .W34TO28(66), .W34TO29(21), .W34TO30(17), .W34TO31(150), .W34TO32(-49), .W34TO33(119), .W34TO34(-189), .W34TO35(130), .W34TO36(-88), .W34TO37(97), .W34TO38(103), .W34TO39(183), .W34TO40(-22), .W34TO41(-45), .W34TO42(108), .W34TO43(70), .W34TO44(157), .W34TO45(112), .W34TO46(134), .W34TO47(49), .W34TO48(54), .W34TO49(-56), .W34TO50(112), .W34TO51(69), .W34TO52(41), .W34TO53(-21), .W34TO54(33), .W34TO55(-63), .W34TO56(16), .W34TO57(-143), .W34TO58(-45), .W34TO59(-44), .W34TO60(51), .W34TO61(-9), .W34TO62(127), .W34TO63(174), .W34TO64(-89), .W34TO65(113), .W34TO66(81), .W34TO67(32), .W34TO68(-95), .W34TO69(179), .W34TO70(-61), .W34TO71(51), .W34TO72(118), .W34TO73(28), .W34TO74(68), .W34TO75(-143), .W34TO76(125), .W34TO77(167), .W34TO78(102), .W34TO79(-154), .W34TO80(-91), .W34TO81(157), .W34TO82(35), .W34TO83(-121), .W34TO84(-28), .W34TO85(124), .W34TO86(106), .W34TO87(-10), .W34TO88(69), .W34TO89(-1), .W34TO90(131), .W34TO91(-1), .W34TO92(-146), .W34TO93(-83), .W34TO94(113), .W34TO95(122), .W34TO96(43), .W34TO97(127), .W34TO98(-49), .W34TO99(99), .W35TO0(51), .W35TO1(-12), .W35TO2(-112), .W35TO3(154), .W35TO4(-146), .W35TO5(117), .W35TO6(-33), .W35TO7(143), .W35TO8(189), .W35TO9(128), .W35TO10(29), .W35TO11(72), .W35TO12(-180), .W35TO13(-34), .W35TO14(150), .W35TO15(139), .W35TO16(18), .W35TO17(56), .W35TO18(-87), .W35TO19(-6), .W35TO20(-192), .W35TO21(-169), .W35TO22(-77), .W35TO23(-186), .W35TO24(133), .W35TO25(-163), .W35TO26(74), .W35TO27(3), .W35TO28(47), .W35TO29(118), .W35TO30(63), .W35TO31(158), .W35TO32(128), .W35TO33(156), .W35TO34(-194), .W35TO35(-17), .W35TO36(165), .W35TO37(-8), .W35TO38(175), .W35TO39(-89), .W35TO40(-211), .W35TO41(58), .W35TO42(-91), .W35TO43(87), .W35TO44(-160), .W35TO45(-36), .W35TO46(23), .W35TO47(80), .W35TO48(-209), .W35TO49(130), .W35TO50(220), .W35TO51(178), .W35TO52(-12), .W35TO53(229), .W35TO54(84), .W35TO55(221), .W35TO56(202), .W35TO57(77), .W35TO58(-87), .W35TO59(18), .W35TO60(151), .W35TO61(17), .W35TO62(122), .W35TO63(-86), .W35TO64(-1), .W35TO65(-25), .W35TO66(-83), .W35TO67(-174), .W35TO68(117), .W35TO69(199), .W35TO70(126), .W35TO71(-17), .W35TO72(-69), .W35TO73(-184), .W35TO74(105), .W35TO75(30), .W35TO76(36), .W35TO77(-104), .W35TO78(-189), .W35TO79(84), .W35TO80(-4), .W35TO81(-87), .W35TO82(-4), .W35TO83(37), .W35TO84(33), .W35TO85(145), .W35TO86(-143), .W35TO87(-5), .W35TO88(165), .W35TO89(84), .W35TO90(-75), .W35TO91(23), .W35TO92(-47), .W35TO93(210), .W35TO94(36), .W35TO95(-59), .W35TO96(-41), .W35TO97(-143), .W35TO98(75), .W35TO99(64), .W36TO0(67), .W36TO1(41), .W36TO2(-173), .W36TO3(-78), .W36TO4(-107), .W36TO5(-91), .W36TO6(-80), .W36TO7(51), .W36TO8(145), .W36TO9(-62), .W36TO10(29), .W36TO11(6), .W36TO12(-90), .W36TO13(-90), .W36TO14(-153), .W36TO15(-64), .W36TO16(120), .W36TO17(107), .W36TO18(125), .W36TO19(115), .W36TO20(18), .W36TO21(13), .W36TO22(-94), .W36TO23(-97), .W36TO24(109), .W36TO25(160), .W36TO26(-86), .W36TO27(57), .W36TO28(164), .W36TO29(-123), .W36TO30(146), .W36TO31(106), .W36TO32(-51), .W36TO33(73), .W36TO34(-97), .W36TO35(136), .W36TO36(26), .W36TO37(43), .W36TO38(111), .W36TO39(21), .W36TO40(-161), .W36TO41(70), .W36TO42(-153), .W36TO43(-40), .W36TO44(56), .W36TO45(144), .W36TO46(-146), .W36TO47(10), .W36TO48(22), .W36TO49(-133), .W36TO50(59), .W36TO51(31), .W36TO52(-181), .W36TO53(11), .W36TO54(-107), .W36TO55(-5), .W36TO56(-115), .W36TO57(-20), .W36TO58(8), .W36TO59(-91), .W36TO60(19), .W36TO61(-14), .W36TO62(-128), .W36TO63(-138), .W36TO64(3), .W36TO65(42), .W36TO66(-214), .W36TO67(-13), .W36TO68(-109), .W36TO69(-141), .W36TO70(89), .W36TO71(-21), .W36TO72(-39), .W36TO73(123), .W36TO74(-29), .W36TO75(-126), .W36TO76(3), .W36TO77(175), .W36TO78(139), .W36TO79(168), .W36TO80(-105), .W36TO81(-5), .W36TO82(-31), .W36TO83(-204), .W36TO84(-19), .W36TO85(10), .W36TO86(147), .W36TO87(-82), .W36TO88(139), .W36TO89(-156), .W36TO90(177), .W36TO91(212), .W36TO92(-18), .W36TO93(200), .W36TO94(-101), .W36TO95(131), .W36TO96(49), .W36TO97(-109), .W36TO98(-123), .W36TO99(-44), .W37TO0(-156), .W37TO1(138), .W37TO2(-191), .W37TO3(-143), .W37TO4(-45), .W37TO5(115), .W37TO6(151), .W37TO7(-65), .W37TO8(-66), .W37TO9(134), .W37TO10(180), .W37TO11(-182), .W37TO12(24), .W37TO13(-94), .W37TO14(158), .W37TO15(160), .W37TO16(205), .W37TO17(-48), .W37TO18(-46), .W37TO19(21), .W37TO20(28), .W37TO21(85), .W37TO22(111), .W37TO23(-140), .W37TO24(-138), .W37TO25(128), .W37TO26(147), .W37TO27(-132), .W37TO28(83), .W37TO29(4), .W37TO30(-16), .W37TO31(12), .W37TO32(192), .W37TO33(41), .W37TO34(-189), .W37TO35(105), .W37TO36(-201), .W37TO37(28), .W37TO38(-60), .W37TO39(64), .W37TO40(-231), .W37TO41(-106), .W37TO42(7), .W37TO43(43), .W37TO44(62), .W37TO45(112), .W37TO46(-145), .W37TO47(-71), .W37TO48(-53), .W37TO49(-70), .W37TO50(140), .W37TO51(218), .W37TO52(-5), .W37TO53(28), .W37TO54(273), .W37TO55(120), .W37TO56(58), .W37TO57(-97), .W37TO58(-161), .W37TO59(33), .W37TO60(94), .W37TO61(-119), .W37TO62(-183), .W37TO63(89), .W37TO64(-177), .W37TO65(-50), .W37TO66(99), .W37TO67(52), .W37TO68(144), .W37TO69(-155), .W37TO70(-161), .W37TO71(-43), .W37TO72(-22), .W37TO73(-102), .W37TO74(-131), .W37TO75(-99), .W37TO76(-93), .W37TO77(77), .W37TO78(-3), .W37TO79(71), .W37TO80(-163), .W37TO81(100), .W37TO82(-147), .W37TO83(52), .W37TO84(140), .W37TO85(-107), .W37TO86(74), .W37TO87(-100), .W37TO88(10), .W37TO89(-82), .W37TO90(114), .W37TO91(206), .W37TO92(-19), .W37TO93(8), .W37TO94(-171), .W37TO95(157), .W37TO96(12), .W37TO97(-35), .W37TO98(-70), .W37TO99(124), .W38TO0(-148), .W38TO1(-51), .W38TO2(-55), .W38TO3(-75), .W38TO4(-79), .W38TO5(32), .W38TO6(-182), .W38TO7(56), .W38TO8(69), .W38TO9(125), .W38TO10(-111), .W38TO11(-116), .W38TO12(114), .W38TO13(41), .W38TO14(21), .W38TO15(158), .W38TO16(-8), .W38TO17(0), .W38TO18(158), .W38TO19(20), .W38TO20(-20), .W38TO21(-58), .W38TO22(-37), .W38TO23(-176), .W38TO24(75), .W38TO25(100), .W38TO26(148), .W38TO27(-95), .W38TO28(-122), .W38TO29(164), .W38TO30(-180), .W38TO31(-85), .W38TO32(134), .W38TO33(84), .W38TO34(-77), .W38TO35(-16), .W38TO36(63), .W38TO37(135), .W38TO38(-53), .W38TO39(-13), .W38TO40(106), .W38TO41(-46), .W38TO42(37), .W38TO43(-83), .W38TO44(183), .W38TO45(54), .W38TO46(59), .W38TO47(-90), .W38TO48(-65), .W38TO49(-97), .W38TO50(-118), .W38TO51(117), .W38TO52(46), .W38TO53(-296), .W38TO54(225), .W38TO55(-54), .W38TO56(-167), .W38TO57(-53), .W38TO58(-94), .W38TO59(197), .W38TO60(103), .W38TO61(20), .W38TO62(63), .W38TO63(-77), .W38TO64(-174), .W38TO65(47), .W38TO66(58), .W38TO67(-152), .W38TO68(-47), .W38TO69(-126), .W38TO70(31), .W38TO71(205), .W38TO72(-160), .W38TO73(14), .W38TO74(-169), .W38TO75(-9), .W38TO76(0), .W38TO77(136), .W38TO78(-76), .W38TO79(-19), .W38TO80(-143), .W38TO81(188), .W38TO82(-63), .W38TO83(40), .W38TO84(-32), .W38TO85(-145), .W38TO86(-86), .W38TO87(3), .W38TO88(2), .W38TO89(128), .W38TO90(-27), .W38TO91(49), .W38TO92(95), .W38TO93(-50), .W38TO94(-49), .W38TO95(36), .W38TO96(-108), .W38TO97(-75), .W38TO98(-121), .W38TO99(153), .W39TO0(-86), .W39TO1(118), .W39TO2(64), .W39TO3(-12), .W39TO4(8), .W39TO5(-170), .W39TO6(137), .W39TO7(-64), .W39TO8(4), .W39TO9(68), .W39TO10(-55), .W39TO11(-180), .W39TO12(-87), .W39TO13(-60), .W39TO14(25), .W39TO15(-128), .W39TO16(-25), .W39TO17(-115), .W39TO18(-80), .W39TO19(64), .W39TO20(138), .W39TO21(-83), .W39TO22(-175), .W39TO23(71), .W39TO24(-161), .W39TO25(-116), .W39TO26(-17), .W39TO27(65), .W39TO28(-119), .W39TO29(-108), .W39TO30(-175), .W39TO31(143), .W39TO32(125), .W39TO33(167), .W39TO34(-154), .W39TO35(-96), .W39TO36(-2), .W39TO37(-82), .W39TO38(-67), .W39TO39(168), .W39TO40(-149), .W39TO41(-108), .W39TO42(-121), .W39TO43(-35), .W39TO44(-65), .W39TO45(59), .W39TO46(-64), .W39TO47(-54), .W39TO48(86), .W39TO49(-68), .W39TO50(134), .W39TO51(48), .W39TO52(142), .W39TO53(-140), .W39TO54(89), .W39TO55(184), .W39TO56(-30), .W39TO57(21), .W39TO58(-39), .W39TO59(58), .W39TO60(1), .W39TO61(-159), .W39TO62(-106), .W39TO63(179), .W39TO64(-35), .W39TO65(149), .W39TO66(4), .W39TO67(-93), .W39TO68(16), .W39TO69(154), .W39TO70(-180), .W39TO71(-68), .W39TO72(-104), .W39TO73(-63), .W39TO74(102), .W39TO75(-36), .W39TO76(75), .W39TO77(163), .W39TO78(-127), .W39TO79(169), .W39TO80(-180), .W39TO81(-73), .W39TO82(177), .W39TO83(74), .W39TO84(-23), .W39TO85(-65), .W39TO86(-180), .W39TO87(187), .W39TO88(-112), .W39TO89(-96), .W39TO90(-70), .W39TO91(65), .W39TO92(66), .W39TO93(174), .W39TO94(101), .W39TO95(-75), .W39TO96(93), .W39TO97(-72), .W39TO98(81), .W39TO99(190), .W40TO0(25), .W40TO1(-24), .W40TO2(-162), .W40TO3(-184), .W40TO4(107), .W40TO5(139), .W40TO6(70), .W40TO7(-134), .W40TO8(9), .W40TO9(-190), .W40TO10(42), .W40TO11(-151), .W40TO12(-32), .W40TO13(-121), .W40TO14(112), .W40TO15(-39), .W40TO16(-65), .W40TO17(144), .W40TO18(173), .W40TO19(63), .W40TO20(98), .W40TO21(-3), .W40TO22(-6), .W40TO23(28), .W40TO24(53), .W40TO25(114), .W40TO26(-73), .W40TO27(-66), .W40TO28(135), .W40TO29(5), .W40TO30(118), .W40TO31(-141), .W40TO32(46), .W40TO33(165), .W40TO34(50), .W40TO35(149), .W40TO36(-99), .W40TO37(179), .W40TO38(168), .W40TO39(31), .W40TO40(-18), .W40TO41(-6), .W40TO42(-171), .W40TO43(180), .W40TO44(26), .W40TO45(119), .W40TO46(-159), .W40TO47(-51), .W40TO48(-60), .W40TO49(-22), .W40TO50(-12), .W40TO51(-82), .W40TO52(-148), .W40TO53(-113), .W40TO54(-178), .W40TO55(-69), .W40TO56(-17), .W40TO57(27), .W40TO58(-188), .W40TO59(-32), .W40TO60(107), .W40TO61(128), .W40TO62(76), .W40TO63(175), .W40TO64(-133), .W40TO65(-134), .W40TO66(-41), .W40TO67(107), .W40TO68(81), .W40TO69(-1), .W40TO70(63), .W40TO71(77), .W40TO72(186), .W40TO73(127), .W40TO74(6), .W40TO75(-96), .W40TO76(51), .W40TO77(165), .W40TO78(-37), .W40TO79(-25), .W40TO80(188), .W40TO81(-181), .W40TO82(-144), .W40TO83(146), .W40TO84(-6), .W40TO85(60), .W40TO86(-155), .W40TO87(98), .W40TO88(99), .W40TO89(-120), .W40TO90(-9), .W40TO91(105), .W40TO92(71), .W40TO93(-182), .W40TO94(65), .W40TO95(53), .W40TO96(-125), .W40TO97(-20), .W40TO98(133), .W40TO99(-39), .W41TO0(124), .W41TO1(-58), .W41TO2(116), .W41TO3(142), .W41TO4(-64), .W41TO5(45), .W41TO6(-157), .W41TO7(69), .W41TO8(-128), .W41TO9(146), .W41TO10(-67), .W41TO11(-107), .W41TO12(-103), .W41TO13(-61), .W41TO14(57), .W41TO15(159), .W41TO16(-130), .W41TO17(-176), .W41TO18(116), .W41TO19(-170), .W41TO20(-79), .W41TO21(-141), .W41TO22(159), .W41TO23(77), .W41TO24(7), .W41TO25(84), .W41TO26(-93), .W41TO27(-108), .W41TO28(111), .W41TO29(137), .W41TO30(-195), .W41TO31(110), .W41TO32(-147), .W41TO33(-198), .W41TO34(-189), .W41TO35(-143), .W41TO36(162), .W41TO37(-141), .W41TO38(30), .W41TO39(112), .W41TO40(19), .W41TO41(132), .W41TO42(-181), .W41TO43(70), .W41TO44(133), .W41TO45(106), .W41TO46(114), .W41TO47(-126), .W41TO48(88), .W41TO49(-60), .W41TO50(181), .W41TO51(208), .W41TO52(-9), .W41TO53(76), .W41TO54(16), .W41TO55(149), .W41TO56(3), .W41TO57(-178), .W41TO58(-146), .W41TO59(136), .W41TO60(-59), .W41TO61(-213), .W41TO62(25), .W41TO63(-220), .W41TO64(-180), .W41TO65(-122), .W41TO66(9), .W41TO67(-94), .W41TO68(-2), .W41TO69(-21), .W41TO70(-178), .W41TO71(-113), .W41TO72(188), .W41TO73(91), .W41TO74(-52), .W41TO75(36), .W41TO76(71), .W41TO77(-38), .W41TO78(100), .W41TO79(21), .W41TO80(-1), .W41TO81(-187), .W41TO82(-18), .W41TO83(-9), .W41TO84(-91), .W41TO85(-15), .W41TO86(-29), .W41TO87(-10), .W41TO88(43), .W41TO89(-176), .W41TO90(-171), .W41TO91(-23), .W41TO92(23), .W41TO93(142), .W41TO94(54), .W41TO95(-8), .W41TO96(-90), .W41TO97(109), .W41TO98(27), .W41TO99(-30), .W42TO0(-118), .W42TO1(1), .W42TO2(126), .W42TO3(154), .W42TO4(200), .W42TO5(-198), .W42TO6(173), .W42TO7(-173), .W42TO8(-12), .W42TO9(146), .W42TO10(164), .W42TO11(127), .W42TO12(-72), .W42TO13(7), .W42TO14(68), .W42TO15(163), .W42TO16(121), .W42TO17(-176), .W42TO18(-110), .W42TO19(-49), .W42TO20(-3), .W42TO21(-55), .W42TO22(8), .W42TO23(91), .W42TO24(-35), .W42TO25(78), .W42TO26(-54), .W42TO27(-8), .W42TO28(-175), .W42TO29(-16), .W42TO30(149), .W42TO31(121), .W42TO32(-54), .W42TO33(140), .W42TO34(-150), .W42TO35(-127), .W42TO36(20), .W42TO37(2), .W42TO38(125), .W42TO39(22), .W42TO40(122), .W42TO41(288), .W42TO42(44), .W42TO43(91), .W42TO44(-98), .W42TO45(-136), .W42TO46(-19), .W42TO47(-100), .W42TO48(-172), .W42TO49(-97), .W42TO50(102), .W42TO51(-54), .W42TO52(140), .W42TO53(58), .W42TO54(29), .W42TO55(136), .W42TO56(32), .W42TO57(-16), .W42TO58(-100), .W42TO59(190), .W42TO60(2), .W42TO61(40), .W42TO62(1), .W42TO63(-42), .W42TO64(-93), .W42TO65(17), .W42TO66(-161), .W42TO67(-76), .W42TO68(210), .W42TO69(-8), .W42TO70(11), .W42TO71(-82), .W42TO72(96), .W42TO73(105), .W42TO74(-101), .W42TO75(155), .W42TO76(118), .W42TO77(-100), .W42TO78(179), .W42TO79(-177), .W42TO80(214), .W42TO81(-26), .W42TO82(-124), .W42TO83(-197), .W42TO84(27), .W42TO85(94), .W42TO86(-216), .W42TO87(34), .W42TO88(-35), .W42TO89(-2), .W42TO90(38), .W42TO91(-109), .W42TO92(205), .W42TO93(36), .W42TO94(-159), .W42TO95(106), .W42TO96(-10), .W42TO97(200), .W42TO98(-6), .W42TO99(31), .W43TO0(-18), .W43TO1(-102), .W43TO2(-140), .W43TO3(126), .W43TO4(6), .W43TO5(-68), .W43TO6(178), .W43TO7(161), .W43TO8(192), .W43TO9(-54), .W43TO10(63), .W43TO11(70), .W43TO12(-66), .W43TO13(-79), .W43TO14(-87), .W43TO15(101), .W43TO16(-107), .W43TO17(119), .W43TO18(-159), .W43TO19(2), .W43TO20(-84), .W43TO21(35), .W43TO22(-83), .W43TO23(-36), .W43TO24(-2), .W43TO25(-53), .W43TO26(-25), .W43TO27(144), .W43TO28(145), .W43TO29(100), .W43TO30(-116), .W43TO31(203), .W43TO32(56), .W43TO33(-119), .W43TO34(-110), .W43TO35(136), .W43TO36(85), .W43TO37(69), .W43TO38(151), .W43TO39(31), .W43TO40(79), .W43TO41(186), .W43TO42(-120), .W43TO43(-120), .W43TO44(52), .W43TO45(-89), .W43TO46(94), .W43TO47(2), .W43TO48(-14), .W43TO49(-306), .W43TO50(24), .W43TO51(-98), .W43TO52(-150), .W43TO53(-12), .W43TO54(2), .W43TO55(31), .W43TO56(87), .W43TO57(-41), .W43TO58(2), .W43TO59(37), .W43TO60(178), .W43TO61(7), .W43TO62(66), .W43TO63(49), .W43TO64(106), .W43TO65(23), .W43TO66(62), .W43TO67(75), .W43TO68(113), .W43TO69(62), .W43TO70(-85), .W43TO71(-263), .W43TO72(163), .W43TO73(-129), .W43TO74(-190), .W43TO75(-96), .W43TO76(-79), .W43TO77(-130), .W43TO78(192), .W43TO79(-128), .W43TO80(43), .W43TO81(-144), .W43TO82(27), .W43TO83(-266), .W43TO84(51), .W43TO85(-20), .W43TO86(-139), .W43TO87(4), .W43TO88(-9), .W43TO89(-48), .W43TO90(135), .W43TO91(-183), .W43TO92(0), .W43TO93(195), .W43TO94(20), .W43TO95(210), .W43TO96(-7), .W43TO97(-107), .W43TO98(95), .W43TO99(76), .W44TO0(-66), .W44TO1(155), .W44TO2(111), .W44TO3(-170), .W44TO4(-231), .W44TO5(-78), .W44TO6(-43), .W44TO7(145), .W44TO8(166), .W44TO9(171), .W44TO10(20), .W44TO11(-3), .W44TO12(173), .W44TO13(-68), .W44TO14(119), .W44TO15(35), .W44TO16(-165), .W44TO17(208), .W44TO18(187), .W44TO19(115), .W44TO20(39), .W44TO21(210), .W44TO22(74), .W44TO23(24), .W44TO24(-36), .W44TO25(-2), .W44TO26(88), .W44TO27(-102), .W44TO28(-126), .W44TO29(-57), .W44TO30(107), .W44TO31(170), .W44TO32(-121), .W44TO33(-62), .W44TO34(149), .W44TO35(170), .W44TO36(140), .W44TO37(59), .W44TO38(81), .W44TO39(-55), .W44TO40(66), .W44TO41(-192), .W44TO42(-173), .W44TO43(-147), .W44TO44(119), .W44TO45(6), .W44TO46(-116), .W44TO47(-36), .W44TO48(-87), .W44TO49(86), .W44TO50(33), .W44TO51(-65), .W44TO52(-202), .W44TO53(-56), .W44TO54(-116), .W44TO55(-5), .W44TO56(190), .W44TO57(-167), .W44TO58(56), .W44TO59(-40), .W44TO60(-40), .W44TO61(136), .W44TO62(-83), .W44TO63(-29), .W44TO64(-71), .W44TO65(-56), .W44TO66(-38), .W44TO67(-59), .W44TO68(13), .W44TO69(-98), .W44TO70(33), .W44TO71(-30), .W44TO72(155), .W44TO73(77), .W44TO74(-32), .W44TO75(-19), .W44TO76(63), .W44TO77(6), .W44TO78(32), .W44TO79(62), .W44TO80(146), .W44TO81(16), .W44TO82(47), .W44TO83(10), .W44TO84(204), .W44TO85(-60), .W44TO86(129), .W44TO87(27), .W44TO88(-137), .W44TO89(-137), .W44TO90(-18), .W44TO91(-103), .W44TO92(-44), .W44TO93(29), .W44TO94(-142), .W44TO95(225), .W44TO96(76), .W44TO97(-222), .W44TO98(13), .W44TO99(-83), .W45TO0(-73), .W45TO1(-79), .W45TO2(-8), .W45TO3(107), .W45TO4(-54), .W45TO5(133), .W45TO6(123), .W45TO7(135), .W45TO8(-30), .W45TO9(-7), .W45TO10(87), .W45TO11(-81), .W45TO12(14), .W45TO13(38), .W45TO14(-155), .W45TO15(148), .W45TO16(10), .W45TO17(-35), .W45TO18(-131), .W45TO19(-89), .W45TO20(-93), .W45TO21(11), .W45TO22(109), .W45TO23(-138), .W45TO24(-11), .W45TO25(228), .W45TO26(88), .W45TO27(-11), .W45TO28(8), .W45TO29(156), .W45TO30(202), .W45TO31(143), .W45TO32(223), .W45TO33(186), .W45TO34(98), .W45TO35(-173), .W45TO36(-127), .W45TO37(-151), .W45TO38(199), .W45TO39(-38), .W45TO40(56), .W45TO41(171), .W45TO42(-75), .W45TO43(-80), .W45TO44(132), .W45TO45(49), .W45TO46(-86), .W45TO47(-89), .W45TO48(-198), .W45TO49(138), .W45TO50(37), .W45TO51(209), .W45TO52(-6), .W45TO53(-33), .W45TO54(-78), .W45TO55(-97), .W45TO56(-131), .W45TO57(-196), .W45TO58(-152), .W45TO59(-55), .W45TO60(-115), .W45TO61(-2), .W45TO62(-37), .W45TO63(58), .W45TO64(-38), .W45TO65(48), .W45TO66(-54), .W45TO67(-76), .W45TO68(150), .W45TO69(29), .W45TO70(85), .W45TO71(96), .W45TO72(147), .W45TO73(21), .W45TO74(60), .W45TO75(9), .W45TO76(81), .W45TO77(20), .W45TO78(-191), .W45TO79(-32), .W45TO80(86), .W45TO81(-52), .W45TO82(69), .W45TO83(-110), .W45TO84(-199), .W45TO85(-17), .W45TO86(79), .W45TO87(202), .W45TO88(-4), .W45TO89(-166), .W45TO90(43), .W45TO91(35), .W45TO92(-116), .W45TO93(180), .W45TO94(96), .W45TO95(-114), .W45TO96(10), .W45TO97(-75), .W45TO98(-185), .W45TO99(97), .W46TO0(59), .W46TO1(130), .W46TO2(106), .W46TO3(-56), .W46TO4(-57), .W46TO5(-28), .W46TO6(62), .W46TO7(-103), .W46TO8(112), .W46TO9(73), .W46TO10(-150), .W46TO11(62), .W46TO12(-77), .W46TO13(128), .W46TO14(148), .W46TO15(33), .W46TO16(-126), .W46TO17(-252), .W46TO18(72), .W46TO19(-132), .W46TO20(64), .W46TO21(-104), .W46TO22(-71), .W46TO23(190), .W46TO24(143), .W46TO25(-150), .W46TO26(-121), .W46TO27(84), .W46TO28(-38), .W46TO29(-73), .W46TO30(157), .W46TO31(-41), .W46TO32(-108), .W46TO33(170), .W46TO34(51), .W46TO35(183), .W46TO36(-52), .W46TO37(-144), .W46TO38(-166), .W46TO39(167), .W46TO40(23), .W46TO41(61), .W46TO42(-165), .W46TO43(108), .W46TO44(104), .W46TO45(26), .W46TO46(-112), .W46TO47(-82), .W46TO48(-110), .W46TO49(182), .W46TO50(14), .W46TO51(-17), .W46TO52(-115), .W46TO53(59), .W46TO54(-20), .W46TO55(153), .W46TO56(94), .W46TO57(-177), .W46TO58(-63), .W46TO59(-47), .W46TO60(-70), .W46TO61(-89), .W46TO62(126), .W46TO63(-49), .W46TO64(102), .W46TO65(-5), .W46TO66(122), .W46TO67(44), .W46TO68(50), .W46TO69(-130), .W46TO70(14), .W46TO71(132), .W46TO72(-21), .W46TO73(-157), .W46TO74(-37), .W46TO75(-41), .W46TO76(80), .W46TO77(-191), .W46TO78(38), .W46TO79(197), .W46TO80(-72), .W46TO81(129), .W46TO82(-96), .W46TO83(-85), .W46TO84(13), .W46TO85(121), .W46TO86(0), .W46TO87(20), .W46TO88(36), .W46TO89(58), .W46TO90(75), .W46TO91(-95), .W46TO92(110), .W46TO93(64), .W46TO94(2), .W46TO95(150), .W46TO96(128), .W46TO97(38), .W46TO98(66), .W46TO99(-137), .W47TO0(-19), .W47TO1(44), .W47TO2(-175), .W47TO3(157), .W47TO4(-150), .W47TO5(170), .W47TO6(146), .W47TO7(89), .W47TO8(180), .W47TO9(27), .W47TO10(28), .W47TO11(-153), .W47TO12(-23), .W47TO13(-162), .W47TO14(62), .W47TO15(-117), .W47TO16(-171), .W47TO17(30), .W47TO18(37), .W47TO19(172), .W47TO20(-171), .W47TO21(-97), .W47TO22(174), .W47TO23(166), .W47TO24(-120), .W47TO25(31), .W47TO26(-68), .W47TO27(-137), .W47TO28(-30), .W47TO29(-4), .W47TO30(54), .W47TO31(109), .W47TO32(54), .W47TO33(95), .W47TO34(76), .W47TO35(40), .W47TO36(81), .W47TO37(90), .W47TO38(-98), .W47TO39(145), .W47TO40(5), .W47TO41(-160), .W47TO42(48), .W47TO43(180), .W47TO44(-12), .W47TO45(190), .W47TO46(-18), .W47TO47(174), .W47TO48(-185), .W47TO49(-24), .W47TO50(184), .W47TO51(147), .W47TO52(52), .W47TO53(-73), .W47TO54(155), .W47TO55(-75), .W47TO56(111), .W47TO57(-52), .W47TO58(53), .W47TO59(19), .W47TO60(-55), .W47TO61(38), .W47TO62(132), .W47TO63(175), .W47TO64(-134), .W47TO65(67), .W47TO66(-159), .W47TO67(-45), .W47TO68(-100), .W47TO69(-168), .W47TO70(-78), .W47TO71(-47), .W47TO72(79), .W47TO73(81), .W47TO74(139), .W47TO75(11), .W47TO76(181), .W47TO77(163), .W47TO78(-175), .W47TO79(-9), .W47TO80(114), .W47TO81(-67), .W47TO82(-31), .W47TO83(-152), .W47TO84(-23), .W47TO85(-65), .W47TO86(44), .W47TO87(-46), .W47TO88(-55), .W47TO89(29), .W47TO90(-105), .W47TO91(188), .W47TO92(105), .W47TO93(144), .W47TO94(102), .W47TO95(163), .W47TO96(-177), .W47TO97(72), .W47TO98(-31), .W47TO99(-179), .W48TO0(35), .W48TO1(183), .W48TO2(-158), .W48TO3(17), .W48TO4(67), .W48TO5(-186), .W48TO6(182), .W48TO7(11), .W48TO8(-35), .W48TO9(-54), .W48TO10(99), .W48TO11(-91), .W48TO12(-128), .W48TO13(106), .W48TO14(-83), .W48TO15(31), .W48TO16(-65), .W48TO17(135), .W48TO18(53), .W48TO19(-88), .W48TO20(-173), .W48TO21(-98), .W48TO22(107), .W48TO23(-63), .W48TO24(149), .W48TO25(-186), .W48TO26(-80), .W48TO27(-128), .W48TO28(-91), .W48TO29(-32), .W48TO30(38), .W48TO31(-97), .W48TO32(-123), .W48TO33(-66), .W48TO34(5), .W48TO35(-123), .W48TO36(53), .W48TO37(-186), .W48TO38(157), .W48TO39(79), .W48TO40(-168), .W48TO41(185), .W48TO42(189), .W48TO43(-69), .W48TO44(-148), .W48TO45(-152), .W48TO46(169), .W48TO47(83), .W48TO48(24), .W48TO49(-139), .W48TO50(-105), .W48TO51(-139), .W48TO52(-136), .W48TO53(171), .W48TO54(182), .W48TO55(117), .W48TO56(9), .W48TO57(122), .W48TO58(-118), .W48TO59(-26), .W48TO60(-10), .W48TO61(180), .W48TO62(168), .W48TO63(-153), .W48TO64(-65), .W48TO65(-59), .W48TO66(-136), .W48TO67(182), .W48TO68(142), .W48TO69(-28), .W48TO70(71), .W48TO71(12), .W48TO72(-88), .W48TO73(-98), .W48TO74(-23), .W48TO75(-23), .W48TO76(35), .W48TO77(-65), .W48TO78(89), .W48TO79(107), .W48TO80(175), .W48TO81(-103), .W48TO82(26), .W48TO83(-28), .W48TO84(-135), .W48TO85(126), .W48TO86(-158), .W48TO87(-98), .W48TO88(42), .W48TO89(34), .W48TO90(157), .W48TO91(153), .W48TO92(117), .W48TO93(-8), .W48TO94(102), .W48TO95(175), .W48TO96(165), .W48TO97(-56), .W48TO98(-46), .W48TO99(-190), .W49TO0(134), .W49TO1(112), .W49TO2(4), .W49TO3(-184), .W49TO4(-184), .W49TO5(121), .W49TO6(-139), .W49TO7(9), .W49TO8(114), .W49TO9(13), .W49TO10(-34), .W49TO11(-182), .W49TO12(37), .W49TO13(122), .W49TO14(147), .W49TO15(137), .W49TO16(-107), .W49TO17(-140), .W49TO18(-104), .W49TO19(-98), .W49TO20(68), .W49TO21(89), .W49TO22(160), .W49TO23(-63), .W49TO24(-94), .W49TO25(183), .W49TO26(110), .W49TO27(-188), .W49TO28(-67), .W49TO29(-116), .W49TO30(146), .W49TO31(28), .W49TO32(111), .W49TO33(-17), .W49TO34(-7), .W49TO35(169), .W49TO36(74), .W49TO37(-6), .W49TO38(-162), .W49TO39(-83), .W49TO40(-137), .W49TO41(129), .W49TO42(185), .W49TO43(87), .W49TO44(186), .W49TO45(-55), .W49TO46(-121), .W49TO47(55), .W49TO48(-74), .W49TO49(-56), .W49TO50(66), .W49TO51(41), .W49TO52(29), .W49TO53(-185), .W49TO54(-66), .W49TO55(75), .W49TO56(-130), .W49TO57(-137), .W49TO58(140), .W49TO59(-133), .W49TO60(-66), .W49TO61(-86), .W49TO62(-170), .W49TO63(106), .W49TO64(157), .W49TO65(-76), .W49TO66(17), .W49TO67(-31), .W49TO68(-136), .W49TO69(141), .W49TO70(129), .W49TO71(161), .W49TO72(-3), .W49TO73(-84), .W49TO74(119), .W49TO75(119), .W49TO76(180), .W49TO77(155), .W49TO78(-1), .W49TO79(168), .W49TO80(174), .W49TO81(-71), .W49TO82(-157), .W49TO83(-152), .W49TO84(115), .W49TO85(67), .W49TO86(-117), .W49TO87(-115), .W49TO88(101), .W49TO89(-140), .W49TO90(-96), .W49TO91(68), .W49TO92(-106), .W49TO93(-89), .W49TO94(-116), .W49TO95(101), .W49TO96(114), .W49TO97(124), .W49TO98(-90), .W49TO99(-48), .W50TO0(-5), .W50TO1(108), .W50TO2(-16), .W50TO3(-26), .W50TO4(-76), .W50TO5(-25), .W50TO6(-36), .W50TO7(29), .W50TO8(-137), .W50TO9(14), .W50TO10(100), .W50TO11(-173), .W50TO12(-52), .W50TO13(31), .W50TO14(149), .W50TO15(-81), .W50TO16(-9), .W50TO17(-22), .W50TO18(-182), .W50TO19(13), .W50TO20(27), .W50TO21(-147), .W50TO22(-166), .W50TO23(-135), .W50TO24(29), .W50TO25(-38), .W50TO26(-139), .W50TO27(20), .W50TO28(-160), .W50TO29(7), .W50TO30(135), .W50TO31(33), .W50TO32(-148), .W50TO33(-130), .W50TO34(6), .W50TO35(66), .W50TO36(135), .W50TO37(206), .W50TO38(207), .W50TO39(-209), .W50TO40(108), .W50TO41(5), .W50TO42(-10), .W50TO43(-57), .W50TO44(-54), .W50TO45(14), .W50TO46(75), .W50TO47(6), .W50TO48(-134), .W50TO49(-101), .W50TO50(-28), .W50TO51(194), .W50TO52(-139), .W50TO53(-164), .W50TO54(65), .W50TO55(-166), .W50TO56(95), .W50TO57(151), .W50TO58(-48), .W50TO59(1), .W50TO60(-151), .W50TO61(197), .W50TO62(-75), .W50TO63(79), .W50TO64(-7), .W50TO65(-189), .W50TO66(34), .W50TO67(101), .W50TO68(-117), .W50TO69(60), .W50TO70(174), .W50TO71(-209), .W50TO72(-56), .W50TO73(-35), .W50TO74(-177), .W50TO75(-49), .W50TO76(-1), .W50TO77(193), .W50TO78(-103), .W50TO79(-137), .W50TO80(203), .W50TO81(118), .W50TO82(27), .W50TO83(-20), .W50TO84(-97), .W50TO85(-160), .W50TO86(-23), .W50TO87(181), .W50TO88(98), .W50TO89(-72), .W50TO90(-138), .W50TO91(7), .W50TO92(-20), .W50TO93(65), .W50TO94(-214), .W50TO95(120), .W50TO96(-93), .W50TO97(4), .W50TO98(125), .W50TO99(115), .W51TO0(-25), .W51TO1(116), .W51TO2(138), .W51TO3(63), .W51TO4(173), .W51TO5(14), .W51TO6(-1), .W51TO7(-45), .W51TO8(112), .W51TO9(42), .W51TO10(49), .W51TO11(166), .W51TO12(-89), .W51TO13(-46), .W51TO14(8), .W51TO15(82), .W51TO16(8), .W51TO17(102), .W51TO18(150), .W51TO19(83), .W51TO20(36), .W51TO21(-8), .W51TO22(-90), .W51TO23(-108), .W51TO24(21), .W51TO25(-161), .W51TO26(-7), .W51TO27(-155), .W51TO28(34), .W51TO29(-186), .W51TO30(135), .W51TO31(-22), .W51TO32(117), .W51TO33(-7), .W51TO34(86), .W51TO35(167), .W51TO36(105), .W51TO37(150), .W51TO38(90), .W51TO39(-98), .W51TO40(-173), .W51TO41(-111), .W51TO42(22), .W51TO43(-28), .W51TO44(43), .W51TO45(98), .W51TO46(128), .W51TO47(-158), .W51TO48(-135), .W51TO49(-259), .W51TO50(-64), .W51TO51(-19), .W51TO52(124), .W51TO53(0), .W51TO54(-92), .W51TO55(52), .W51TO56(25), .W51TO57(-147), .W51TO58(168), .W51TO59(173), .W51TO60(11), .W51TO61(-146), .W51TO62(-193), .W51TO63(147), .W51TO64(173), .W51TO65(-152), .W51TO66(-155), .W51TO67(34), .W51TO68(199), .W51TO69(-101), .W51TO70(0), .W51TO71(13), .W51TO72(102), .W51TO73(-104), .W51TO74(-107), .W51TO75(90), .W51TO76(-154), .W51TO77(-39), .W51TO78(39), .W51TO79(-157), .W51TO80(12), .W51TO81(8), .W51TO82(-27), .W51TO83(78), .W51TO84(-151), .W51TO85(-20), .W51TO86(54), .W51TO87(-84), .W51TO88(110), .W51TO89(160), .W51TO90(189), .W51TO91(-89), .W51TO92(106), .W51TO93(129), .W51TO94(-87), .W51TO95(84), .W51TO96(145), .W51TO97(-32), .W51TO98(-23), .W51TO99(145), .W52TO0(-6), .W52TO1(192), .W52TO2(131), .W52TO3(4), .W52TO4(11), .W52TO5(-51), .W52TO6(-12), .W52TO7(-139), .W52TO8(-111), .W52TO9(-52), .W52TO10(72), .W52TO11(27), .W52TO12(11), .W52TO13(-3), .W52TO14(140), .W52TO15(52), .W52TO16(-41), .W52TO17(-7), .W52TO18(174), .W52TO19(-101), .W52TO20(-13), .W52TO21(-80), .W52TO22(-121), .W52TO23(-55), .W52TO24(75), .W52TO25(-134), .W52TO26(0), .W52TO27(58), .W52TO28(-13), .W52TO29(95), .W52TO30(-73), .W52TO31(81), .W52TO32(-70), .W52TO33(-83), .W52TO34(-90), .W52TO35(10), .W52TO36(142), .W52TO37(-35), .W52TO38(198), .W52TO39(-8), .W52TO40(47), .W52TO41(9), .W52TO42(86), .W52TO43(234), .W52TO44(67), .W52TO45(64), .W52TO46(-88), .W52TO47(-227), .W52TO48(124), .W52TO49(46), .W52TO50(-46), .W52TO51(-6), .W52TO52(-33), .W52TO53(62), .W52TO54(-157), .W52TO55(-107), .W52TO56(-12), .W52TO57(110), .W52TO58(117), .W52TO59(-12), .W52TO60(9), .W52TO61(-91), .W52TO62(46), .W52TO63(-55), .W52TO64(54), .W52TO65(148), .W52TO66(-19), .W52TO67(249), .W52TO68(-131), .W52TO69(24), .W52TO70(-132), .W52TO71(49), .W52TO72(-80), .W52TO73(56), .W52TO74(97), .W52TO75(101), .W52TO76(205), .W52TO77(-20), .W52TO78(148), .W52TO79(-112), .W52TO80(-4), .W52TO81(-16), .W52TO82(65), .W52TO83(113), .W52TO84(-57), .W52TO85(-10), .W52TO86(-67), .W52TO87(-64), .W52TO88(-153), .W52TO89(63), .W52TO90(26), .W52TO91(-80), .W52TO92(194), .W52TO93(-42), .W52TO94(45), .W52TO95(142), .W52TO96(-10), .W52TO97(-81), .W52TO98(-5), .W52TO99(93), .W53TO0(-168), .W53TO1(75), .W53TO2(-25), .W53TO3(-140), .W53TO4(217), .W53TO5(-154), .W53TO6(126), .W53TO7(-227), .W53TO8(-125), .W53TO9(-4), .W53TO10(43), .W53TO11(-42), .W53TO12(36), .W53TO13(129), .W53TO14(-83), .W53TO15(9), .W53TO16(-167), .W53TO17(-91), .W53TO18(-41), .W53TO19(260), .W53TO20(73), .W53TO21(58), .W53TO22(55), .W53TO23(153), .W53TO24(-75), .W53TO25(-110), .W53TO26(-133), .W53TO27(10), .W53TO28(-88), .W53TO29(-183), .W53TO30(-84), .W53TO31(-160), .W53TO32(167), .W53TO33(-61), .W53TO34(-44), .W53TO35(169), .W53TO36(-136), .W53TO37(71), .W53TO38(-136), .W53TO39(-171), .W53TO40(-54), .W53TO41(212), .W53TO42(61), .W53TO43(-93), .W53TO44(-66), .W53TO45(-107), .W53TO46(-13), .W53TO47(69), .W53TO48(97), .W53TO49(71), .W53TO50(-139), .W53TO51(139), .W53TO52(-70), .W53TO53(175), .W53TO54(191), .W53TO55(-68), .W53TO56(91), .W53TO57(-119), .W53TO58(35), .W53TO59(166), .W53TO60(-14), .W53TO61(1), .W53TO62(-67), .W53TO63(-94), .W53TO64(125), .W53TO65(-61), .W53TO66(-197), .W53TO67(180), .W53TO68(-50), .W53TO69(164), .W53TO70(64), .W53TO71(132), .W53TO72(91), .W53TO73(-110), .W53TO74(-1), .W53TO75(-73), .W53TO76(154), .W53TO77(-115), .W53TO78(109), .W53TO79(-23), .W53TO80(4), .W53TO81(-126), .W53TO82(193), .W53TO83(15), .W53TO84(4), .W53TO85(-126), .W53TO86(-81), .W53TO87(-31), .W53TO88(82), .W53TO89(209), .W53TO90(127), .W53TO91(27), .W53TO92(100), .W53TO93(-35), .W53TO94(-127), .W53TO95(135), .W53TO96(-36), .W53TO97(-137), .W53TO98(203), .W53TO99(-181), .W54TO0(124), .W54TO1(-54), .W54TO2(141), .W54TO3(135), .W54TO4(153), .W54TO5(68), .W54TO6(-161), .W54TO7(115), .W54TO8(-178), .W54TO9(-76), .W54TO10(-155), .W54TO11(79), .W54TO12(-156), .W54TO13(-57), .W54TO14(-151), .W54TO15(-31), .W54TO16(99), .W54TO17(32), .W54TO18(144), .W54TO19(149), .W54TO20(-70), .W54TO21(-44), .W54TO22(63), .W54TO23(121), .W54TO24(-4), .W54TO25(19), .W54TO26(92), .W54TO27(165), .W54TO28(-9), .W54TO29(121), .W54TO30(-94), .W54TO31(121), .W54TO32(-104), .W54TO33(-44), .W54TO34(152), .W54TO35(145), .W54TO36(53), .W54TO37(-48), .W54TO38(-33), .W54TO39(-126), .W54TO40(69), .W54TO41(-69), .W54TO42(88), .W54TO43(59), .W54TO44(98), .W54TO45(-106), .W54TO46(37), .W54TO47(-91), .W54TO48(136), .W54TO49(-111), .W54TO50(13), .W54TO51(52), .W54TO52(81), .W54TO53(106), .W54TO54(-17), .W54TO55(1), .W54TO56(165), .W54TO57(78), .W54TO58(9), .W54TO59(141), .W54TO60(9), .W54TO61(-63), .W54TO62(-177), .W54TO63(157), .W54TO64(69), .W54TO65(-137), .W54TO66(66), .W54TO67(84), .W54TO68(126), .W54TO69(79), .W54TO70(118), .W54TO71(131), .W54TO72(159), .W54TO73(11), .W54TO74(-105), .W54TO75(129), .W54TO76(27), .W54TO77(68), .W54TO78(-117), .W54TO79(-74), .W54TO80(-89), .W54TO81(51), .W54TO82(27), .W54TO83(61), .W54TO84(-157), .W54TO85(35), .W54TO86(178), .W54TO87(104), .W54TO88(-13), .W54TO89(211), .W54TO90(-38), .W54TO91(-14), .W54TO92(-64), .W54TO93(-139), .W54TO94(50), .W54TO95(-135), .W54TO96(-76), .W54TO97(20), .W54TO98(-126), .W54TO99(125), .W55TO0(93), .W55TO1(-46), .W55TO2(167), .W55TO3(-123), .W55TO4(113), .W55TO5(-144), .W55TO6(-181), .W55TO7(-79), .W55TO8(25), .W55TO9(-4), .W55TO10(-147), .W55TO11(-62), .W55TO12(42), .W55TO13(-32), .W55TO14(-177), .W55TO15(-180), .W55TO16(-175), .W55TO17(132), .W55TO18(171), .W55TO19(176), .W55TO20(49), .W55TO21(-68), .W55TO22(146), .W55TO23(23), .W55TO24(-27), .W55TO25(15), .W55TO26(100), .W55TO27(-114), .W55TO28(-36), .W55TO29(157), .W55TO30(-166), .W55TO31(164), .W55TO32(-53), .W55TO33(-173), .W55TO34(-98), .W55TO35(-54), .W55TO36(98), .W55TO37(-98), .W55TO38(-56), .W55TO39(115), .W55TO40(-20), .W55TO41(40), .W55TO42(176), .W55TO43(-76), .W55TO44(162), .W55TO45(29), .W55TO46(-34), .W55TO47(-15), .W55TO48(37), .W55TO49(-188), .W55TO50(38), .W55TO51(126), .W55TO52(-84), .W55TO53(159), .W55TO54(163), .W55TO55(92), .W55TO56(37), .W55TO57(-79), .W55TO58(60), .W55TO59(173), .W55TO60(115), .W55TO61(121), .W55TO62(-114), .W55TO63(-45), .W55TO64(92), .W55TO65(7), .W55TO66(-136), .W55TO67(-13), .W55TO68(40), .W55TO69(-83), .W55TO70(178), .W55TO71(50), .W55TO72(189), .W55TO73(83), .W55TO74(-116), .W55TO75(-101), .W55TO76(-33), .W55TO77(125), .W55TO78(52), .W55TO79(99), .W55TO80(-61), .W55TO81(142), .W55TO82(-91), .W55TO83(2), .W55TO84(43), .W55TO85(-4), .W55TO86(108), .W55TO87(-32), .W55TO88(156), .W55TO89(-25), .W55TO90(-122), .W55TO91(-150), .W55TO92(41), .W55TO93(-158), .W55TO94(160), .W55TO95(53), .W55TO96(119), .W55TO97(-131), .W55TO98(-52), .W55TO99(-13), .W56TO0(16), .W56TO1(64), .W56TO2(-119), .W56TO3(-87), .W56TO4(135), .W56TO5(31), .W56TO6(-11), .W56TO7(3), .W56TO8(-186), .W56TO9(-101), .W56TO10(42), .W56TO11(-10), .W56TO12(-78), .W56TO13(108), .W56TO14(-121), .W56TO15(-22), .W56TO16(19), .W56TO17(-100), .W56TO18(-89), .W56TO19(185), .W56TO20(-37), .W56TO21(-118), .W56TO22(-165), .W56TO23(-174), .W56TO24(147), .W56TO25(-20), .W56TO26(-90), .W56TO27(38), .W56TO28(-138), .W56TO29(-1), .W56TO30(45), .W56TO31(-3), .W56TO32(-99), .W56TO33(-64), .W56TO34(-56), .W56TO35(66), .W56TO36(-189), .W56TO37(31), .W56TO38(160), .W56TO39(63), .W56TO40(110), .W56TO41(-124), .W56TO42(-76), .W56TO43(-21), .W56TO44(165), .W56TO45(-110), .W56TO46(-53), .W56TO47(57), .W56TO48(133), .W56TO49(-43), .W56TO50(26), .W56TO51(118), .W56TO52(127), .W56TO53(-123), .W56TO54(171), .W56TO55(-124), .W56TO56(-135), .W56TO57(104), .W56TO58(-60), .W56TO59(-46), .W56TO60(79), .W56TO61(116), .W56TO62(-28), .W56TO63(-161), .W56TO64(38), .W56TO65(158), .W56TO66(70), .W56TO67(-141), .W56TO68(98), .W56TO69(-160), .W56TO70(-188), .W56TO71(-120), .W56TO72(-114), .W56TO73(-149), .W56TO74(134), .W56TO75(-43), .W56TO76(-132), .W56TO77(-30), .W56TO78(-34), .W56TO79(73), .W56TO80(-72), .W56TO81(-15), .W56TO82(-85), .W56TO83(137), .W56TO84(-105), .W56TO85(25), .W56TO86(13), .W56TO87(185), .W56TO88(100), .W56TO89(-130), .W56TO90(77), .W56TO91(-56), .W56TO92(1), .W56TO93(-27), .W56TO94(-176), .W56TO95(8), .W56TO96(-52), .W56TO97(-32), .W56TO98(172), .W56TO99(1), .W57TO0(-75), .W57TO1(7), .W57TO2(93), .W57TO3(-39), .W57TO4(-117), .W57TO5(23), .W57TO6(-129), .W57TO7(176), .W57TO8(-128), .W57TO9(172), .W57TO10(59), .W57TO11(-61), .W57TO12(-8), .W57TO13(-97), .W57TO14(-165), .W57TO15(-124), .W57TO16(-122), .W57TO17(-154), .W57TO18(-144), .W57TO19(-17), .W57TO20(126), .W57TO21(-72), .W57TO22(-65), .W57TO23(163), .W57TO24(-69), .W57TO25(105), .W57TO26(-58), .W57TO27(-53), .W57TO28(-180), .W57TO29(83), .W57TO30(-100), .W57TO31(129), .W57TO32(-27), .W57TO33(94), .W57TO34(-132), .W57TO35(-98), .W57TO36(-101), .W57TO37(78), .W57TO38(34), .W57TO39(-151), .W57TO40(102), .W57TO41(-92), .W57TO42(16), .W57TO43(35), .W57TO44(-92), .W57TO45(-21), .W57TO46(156), .W57TO47(39), .W57TO48(-82), .W57TO49(74), .W57TO50(0), .W57TO51(146), .W57TO52(33), .W57TO53(-156), .W57TO54(40), .W57TO55(-13), .W57TO56(-11), .W57TO57(-93), .W57TO58(-111), .W57TO59(152), .W57TO60(-163), .W57TO61(64), .W57TO62(120), .W57TO63(-100), .W57TO64(150), .W57TO65(129), .W57TO66(-66), .W57TO67(116), .W57TO68(35), .W57TO69(188), .W57TO70(181), .W57TO71(-69), .W57TO72(37), .W57TO73(-154), .W57TO74(-182), .W57TO75(-118), .W57TO76(187), .W57TO77(44), .W57TO78(122), .W57TO79(-46), .W57TO80(12), .W57TO81(77), .W57TO82(127), .W57TO83(110), .W57TO84(-86), .W57TO85(99), .W57TO86(-48), .W57TO87(-121), .W57TO88(-22), .W57TO89(-143), .W57TO90(-151), .W57TO91(143), .W57TO92(-113), .W57TO93(-164), .W57TO94(-62), .W57TO95(-163), .W57TO96(-73), .W57TO97(-56), .W57TO98(-68), .W57TO99(128), .W58TO0(-31), .W58TO1(-133), .W58TO2(-135), .W58TO3(26), .W58TO4(124), .W58TO5(207), .W58TO6(-156), .W58TO7(-59), .W58TO8(21), .W58TO9(186), .W58TO10(189), .W58TO11(134), .W58TO12(-39), .W58TO13(-39), .W58TO14(174), .W58TO15(-8), .W58TO16(30), .W58TO17(-76), .W58TO18(37), .W58TO19(139), .W58TO20(117), .W58TO21(-152), .W58TO22(69), .W58TO23(-196), .W58TO24(224), .W58TO25(49), .W58TO26(-21), .W58TO27(-32), .W58TO28(-30), .W58TO29(-43), .W58TO30(-140), .W58TO31(-207), .W58TO32(117), .W58TO33(28), .W58TO34(21), .W58TO35(-8), .W58TO36(21), .W58TO37(-120), .W58TO38(-128), .W58TO39(112), .W58TO40(-190), .W58TO41(-38), .W58TO42(-155), .W58TO43(-48), .W58TO44(-98), .W58TO45(-35), .W58TO46(92), .W58TO47(24), .W58TO48(-167), .W58TO49(-16), .W58TO50(117), .W58TO51(176), .W58TO52(-58), .W58TO53(41), .W58TO54(-78), .W58TO55(-58), .W58TO56(152), .W58TO57(-149), .W58TO58(-123), .W58TO59(45), .W58TO60(48), .W58TO61(-86), .W58TO62(-172), .W58TO63(32), .W58TO64(-90), .W58TO65(-100), .W58TO66(-57), .W58TO67(9), .W58TO68(29), .W58TO69(-152), .W58TO70(-122), .W58TO71(-197), .W58TO72(-95), .W58TO73(130), .W58TO74(-172), .W58TO75(114), .W58TO76(84), .W58TO77(123), .W58TO78(39), .W58TO79(185), .W58TO80(-145), .W58TO81(181), .W58TO82(97), .W58TO83(172), .W58TO84(-101), .W58TO85(-174), .W58TO86(-150), .W58TO87(-9), .W58TO88(-97), .W58TO89(214), .W58TO90(-11), .W58TO91(29), .W58TO92(-119), .W58TO93(12), .W58TO94(57), .W58TO95(-11), .W58TO96(-152), .W58TO97(112), .W58TO98(-119), .W58TO99(170), .W59TO0(148), .W59TO1(-168), .W59TO2(-34), .W59TO3(-104), .W59TO4(-83), .W59TO5(43), .W59TO6(149), .W59TO7(-204), .W59TO8(-16), .W59TO9(16), .W59TO10(25), .W59TO11(16), .W59TO12(174), .W59TO13(126), .W59TO14(159), .W59TO15(-46), .W59TO16(-81), .W59TO17(8), .W59TO18(-37), .W59TO19(9), .W59TO20(113), .W59TO21(61), .W59TO22(86), .W59TO23(36), .W59TO24(152), .W59TO25(-146), .W59TO26(-111), .W59TO27(-92), .W59TO28(132), .W59TO29(50), .W59TO30(-133), .W59TO31(147), .W59TO32(7), .W59TO33(-21), .W59TO34(-200), .W59TO35(72), .W59TO36(-92), .W59TO37(205), .W59TO38(-29), .W59TO39(-208), .W59TO40(-149), .W59TO41(-35), .W59TO42(-172), .W59TO43(155), .W59TO44(92), .W59TO45(-196), .W59TO46(-125), .W59TO47(95), .W59TO48(-121), .W59TO49(145), .W59TO50(9), .W59TO51(70), .W59TO52(26), .W59TO53(-29), .W59TO54(-170), .W59TO55(-174), .W59TO56(67), .W59TO57(144), .W59TO58(-87), .W59TO59(-93), .W59TO60(-142), .W59TO61(-32), .W59TO62(73), .W59TO63(74), .W59TO64(-44), .W59TO65(-177), .W59TO66(-65), .W59TO67(38), .W59TO68(0), .W59TO69(80), .W59TO70(93), .W59TO71(65), .W59TO72(26), .W59TO73(101), .W59TO74(110), .W59TO75(-165), .W59TO76(-47), .W59TO77(-62), .W59TO78(14), .W59TO79(-130), .W59TO80(-85), .W59TO81(-29), .W59TO82(36), .W59TO83(1), .W59TO84(14), .W59TO85(42), .W59TO86(-93), .W59TO87(17), .W59TO88(-41), .W59TO89(226), .W59TO90(51), .W59TO91(-31), .W59TO92(-10), .W59TO93(80), .W59TO94(100), .W59TO95(-191), .W59TO96(-186), .W59TO97(29), .W59TO98(-87), .W59TO99(-13), .W60TO0(-176), .W60TO1(33), .W60TO2(-88), .W60TO3(-230), .W60TO4(-4), .W60TO5(-36), .W60TO6(69), .W60TO7(-172), .W60TO8(55), .W60TO9(-23), .W60TO10(181), .W60TO11(176), .W60TO12(-117), .W60TO13(-50), .W60TO14(-157), .W60TO15(-165), .W60TO16(24), .W60TO17(-134), .W60TO18(147), .W60TO19(201), .W60TO20(75), .W60TO21(-31), .W60TO22(-196), .W60TO23(62), .W60TO24(-78), .W60TO25(-110), .W60TO26(-211), .W60TO27(-125), .W60TO28(-142), .W60TO29(-136), .W60TO30(-97), .W60TO31(-150), .W60TO32(118), .W60TO33(68), .W60TO34(-25), .W60TO35(-41), .W60TO36(19), .W60TO37(-120), .W60TO38(76), .W60TO39(49), .W60TO40(51), .W60TO41(51), .W60TO42(-237), .W60TO43(250), .W60TO44(183), .W60TO45(20), .W60TO46(-47), .W60TO47(-54), .W60TO48(-134), .W60TO49(45), .W60TO50(-105), .W60TO51(-73), .W60TO52(181), .W60TO53(142), .W60TO54(2), .W60TO55(-47), .W60TO56(162), .W60TO57(-108), .W60TO58(-164), .W60TO59(-33), .W60TO60(-40), .W60TO61(-72), .W60TO62(-85), .W60TO63(-44), .W60TO64(-82), .W60TO65(-62), .W60TO66(-199), .W60TO67(137), .W60TO68(-29), .W60TO69(-14), .W60TO70(98), .W60TO71(-106), .W60TO72(208), .W60TO73(-131), .W60TO74(-116), .W60TO75(-186), .W60TO76(-90), .W60TO77(4), .W60TO78(-166), .W60TO79(-52), .W60TO80(46), .W60TO81(51), .W60TO82(54), .W60TO83(-7), .W60TO84(-143), .W60TO85(52), .W60TO86(208), .W60TO87(-96), .W60TO88(135), .W60TO89(-29), .W60TO90(67), .W60TO91(166), .W60TO92(196), .W60TO93(123), .W60TO94(-220), .W60TO95(20), .W60TO96(77), .W60TO97(-63), .W60TO98(204), .W60TO99(85), .W61TO0(-142), .W61TO1(157), .W61TO2(27), .W61TO3(-194), .W61TO4(-70), .W61TO5(-31), .W61TO6(-58), .W61TO7(-132), .W61TO8(-68), .W61TO9(82), .W61TO10(-55), .W61TO11(-142), .W61TO12(-173), .W61TO13(-15), .W61TO14(-94), .W61TO15(186), .W61TO16(97), .W61TO17(-110), .W61TO18(1), .W61TO19(35), .W61TO20(-89), .W61TO21(-69), .W61TO22(95), .W61TO23(129), .W61TO24(11), .W61TO25(241), .W61TO26(158), .W61TO27(-187), .W61TO28(-80), .W61TO29(-151), .W61TO30(187), .W61TO31(47), .W61TO32(200), .W61TO33(-86), .W61TO34(-25), .W61TO35(-151), .W61TO36(32), .W61TO37(125), .W61TO38(-54), .W61TO39(-207), .W61TO40(-114), .W61TO41(6), .W61TO42(-149), .W61TO43(123), .W61TO44(107), .W61TO45(-83), .W61TO46(-2), .W61TO47(30), .W61TO48(-25), .W61TO49(4), .W61TO50(-69), .W61TO51(-1), .W61TO52(198), .W61TO53(-39), .W61TO54(26), .W61TO55(-2), .W61TO56(145), .W61TO57(153), .W61TO58(195), .W61TO59(-102), .W61TO60(-45), .W61TO61(97), .W61TO62(56), .W61TO63(64), .W61TO64(-127), .W61TO65(-31), .W61TO66(-116), .W61TO67(179), .W61TO68(-8), .W61TO69(41), .W61TO70(35), .W61TO71(-99), .W61TO72(199), .W61TO73(34), .W61TO74(170), .W61TO75(-92), .W61TO76(122), .W61TO77(-105), .W61TO78(170), .W61TO79(-4), .W61TO80(86), .W61TO81(-80), .W61TO82(238), .W61TO83(93), .W61TO84(138), .W61TO85(140), .W61TO86(-90), .W61TO87(-211), .W61TO88(-16), .W61TO89(112), .W61TO90(-23), .W61TO91(115), .W61TO92(-70), .W61TO93(-30), .W61TO94(87), .W61TO95(99), .W61TO96(0), .W61TO97(-103), .W61TO98(159), .W61TO99(105), .W62TO0(-59), .W62TO1(-10), .W62TO2(-130), .W62TO3(167), .W62TO4(156), .W62TO5(-214), .W62TO6(39), .W62TO7(116), .W62TO8(-156), .W62TO9(-45), .W62TO10(-80), .W62TO11(-64), .W62TO12(115), .W62TO13(195), .W62TO14(2), .W62TO15(136), .W62TO16(-94), .W62TO17(111), .W62TO18(187), .W62TO19(106), .W62TO20(-179), .W62TO21(-145), .W62TO22(-163), .W62TO23(113), .W62TO24(80), .W62TO25(197), .W62TO26(33), .W62TO27(0), .W62TO28(-152), .W62TO29(-51), .W62TO30(-193), .W62TO31(129), .W62TO32(168), .W62TO33(-51), .W62TO34(96), .W62TO35(37), .W62TO36(-38), .W62TO37(160), .W62TO38(148), .W62TO39(163), .W62TO40(-126), .W62TO41(1), .W62TO42(28), .W62TO43(-75), .W62TO44(60), .W62TO45(-70), .W62TO46(-163), .W62TO47(-33), .W62TO48(-14), .W62TO49(119), .W62TO50(159), .W62TO51(-22), .W62TO52(40), .W62TO53(97), .W62TO54(4), .W62TO55(223), .W62TO56(-160), .W62TO57(103), .W62TO58(-52), .W62TO59(71), .W62TO60(112), .W62TO61(-139), .W62TO62(-144), .W62TO63(-25), .W62TO64(-183), .W62TO65(17), .W62TO66(72), .W62TO67(211), .W62TO68(-130), .W62TO69(68), .W62TO70(214), .W62TO71(104), .W62TO72(67), .W62TO73(-46), .W62TO74(-179), .W62TO75(-40), .W62TO76(212), .W62TO77(-181), .W62TO78(94), .W62TO79(-92), .W62TO80(63), .W62TO81(-83), .W62TO82(207), .W62TO83(-111), .W62TO84(41), .W62TO85(24), .W62TO86(-44), .W62TO87(-113), .W62TO88(134), .W62TO89(-116), .W62TO90(-104), .W62TO91(-138), .W62TO92(-94), .W62TO93(95), .W62TO94(133), .W62TO95(-23), .W62TO96(-118), .W62TO97(-22), .W62TO98(96), .W62TO99(49), .W63TO0(-26), .W63TO1(-128), .W63TO2(216), .W63TO3(24), .W63TO4(-30), .W63TO5(-182), .W63TO6(16), .W63TO7(14), .W63TO8(133), .W63TO9(187), .W63TO10(97), .W63TO11(-81), .W63TO12(-138), .W63TO13(139), .W63TO14(-147), .W63TO15(-87), .W63TO16(-183), .W63TO17(-64), .W63TO18(-96), .W63TO19(70), .W63TO20(161), .W63TO21(-75), .W63TO22(-73), .W63TO23(-17), .W63TO24(2), .W63TO25(34), .W63TO26(127), .W63TO27(3), .W63TO28(104), .W63TO29(-144), .W63TO30(72), .W63TO31(-122), .W63TO32(-102), .W63TO33(-50), .W63TO34(-71), .W63TO35(49), .W63TO36(-131), .W63TO37(-149), .W63TO38(-78), .W63TO39(19), .W63TO40(-140), .W63TO41(27), .W63TO42(143), .W63TO43(135), .W63TO44(-168), .W63TO45(150), .W63TO46(32), .W63TO47(102), .W63TO48(-85), .W63TO49(-121), .W63TO50(188), .W63TO51(10), .W63TO52(-144), .W63TO53(17), .W63TO54(-139), .W63TO55(-104), .W63TO56(169), .W63TO57(140), .W63TO58(123), .W63TO59(145), .W63TO60(143), .W63TO61(-146), .W63TO62(53), .W63TO63(91), .W63TO64(-62), .W63TO65(-123), .W63TO66(-51), .W63TO67(83), .W63TO68(140), .W63TO69(65), .W63TO70(99), .W63TO71(87), .W63TO72(137), .W63TO73(89), .W63TO74(157), .W63TO75(-139), .W63TO76(-154), .W63TO77(-160), .W63TO78(140), .W63TO79(50), .W63TO80(-27), .W63TO81(-153), .W63TO82(57), .W63TO83(-46), .W63TO84(38), .W63TO85(-111), .W63TO86(-128), .W63TO87(-75), .W63TO88(5), .W63TO89(-163), .W63TO90(2), .W63TO91(-182), .W63TO92(115), .W63TO93(-166), .W63TO94(70), .W63TO95(-50), .W63TO96(-89), .W63TO97(-126), .W63TO98(-84), .W63TO99(-4)) layer0(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out0(con0[0]), .out1(con0[1]), .out2(con0[2]), .out3(con0[3]), .out4(con0[4]), .out5(con0[5]), .out6(con0[6]), .out7(con0[7]), .out8(con0[8]), .out9(con0[9]), .out10(con0[10]), .out11(con0[11]), .out12(con0[12]), .out13(con0[13]), .out14(con0[14]), .out15(con0[15]), .out16(con0[16]), .out17(con0[17]), .out18(con0[18]), .out19(con0[19]), .out20(con0[20]), .out21(con0[21]), .out22(con0[22]), .out23(con0[23]), .out24(con0[24]), .out25(con0[25]), .out26(con0[26]), .out27(con0[27]), .out28(con0[28]), .out29(con0[29]), .out30(con0[30]), .out31(con0[31]), .out32(con0[32]), .out33(con0[33]), .out34(con0[34]), .out35(con0[35]), .out36(con0[36]), .out37(con0[37]), .out38(con0[38]), .out39(con0[39]), .out40(con0[40]), .out41(con0[41]), .out42(con0[42]), .out43(con0[43]), .out44(con0[44]), .out45(con0[45]), .out46(con0[46]), .out47(con0[47]), .out48(con0[48]), .out49(con0[49]), .out50(con0[50]), .out51(con0[51]), .out52(con0[52]), .out53(con0[53]), .out54(con0[54]), .out55(con0[55]), .out56(con0[56]), .out57(con0[57]), .out58(con0[58]), .out59(con0[59]), .out60(con0[60]), .out61(con0[61]), .out62(con0[62]), .out63(con0[63]), .out64(con0[64]), .out65(con0[65]), .out66(con0[66]), .out67(con0[67]), .out68(con0[68]), .out69(con0[69]), .out70(con0[70]), .out71(con0[71]), .out72(con0[72]), .out73(con0[73]), .out74(con0[74]), .out75(con0[75]), .out76(con0[76]), .out77(con0[77]), .out78(con0[78]), .out79(con0[79]), .out80(con0[80]), .out81(con0[81]), .out82(con0[82]), .out83(con0[83]), .out84(con0[84]), .out85(con0[85]), .out86(con0[86]), .out87(con0[87]), .out88(con0[88]), .out89(con0[89]), .out90(con0[90]), .out91(con0[91]), .out92(con0[92]), .out93(con0[93]), .out94(con0[94]), .out95(con0[95]), .out96(con0[96]), .out97(con0[97]), .out98(con0[98]), .out99(con0[99]));
layer100in10out #(.W0TO0(261), .W0TO1(214), .W0TO2(256), .W0TO3(263), .W0TO4(66), .W0TO5(-70), .W0TO6(114), .W0TO7(-142), .W0TO8(299), .W0TO9(69), .W1TO0(-113), .W1TO1(-148), .W1TO2(-6), .W1TO3(60), .W1TO4(-146), .W1TO5(-30), .W1TO6(-178), .W1TO7(-85), .W1TO8(120), .W1TO9(-125), .W2TO0(377), .W2TO1(80), .W2TO2(300), .W2TO3(-127), .W2TO4(-205), .W2TO5(-68), .W2TO6(-40), .W2TO7(-72), .W2TO8(5), .W2TO9(-121), .W3TO0(-167), .W3TO1(94), .W3TO2(16), .W3TO3(167), .W3TO4(142), .W3TO5(80), .W3TO6(227), .W3TO7(50), .W3TO8(-21), .W3TO9(195), .W4TO0(170), .W4TO1(178), .W4TO2(300), .W4TO3(-170), .W4TO4(-27), .W4TO5(-218), .W4TO6(359), .W4TO7(-103), .W4TO8(-94), .W4TO9(176), .W5TO0(11), .W5TO1(-163), .W5TO2(7), .W5TO3(-16), .W5TO4(113), .W5TO5(469), .W5TO6(-69), .W5TO7(-147), .W5TO8(-73), .W5TO9(-223), .W6TO0(-81), .W6TO1(-277), .W6TO2(-142), .W6TO3(-24), .W6TO4(-155), .W6TO5(-218), .W6TO6(-148), .W6TO7(-164), .W6TO8(159), .W6TO9(42), .W7TO0(150), .W7TO1(-48), .W7TO2(-18), .W7TO3(112), .W7TO4(-264), .W7TO5(47), .W7TO6(-100), .W7TO7(514), .W7TO8(-233), .W7TO9(5), .W8TO0(-58), .W8TO1(-153), .W8TO2(-90), .W8TO3(-230), .W8TO4(81), .W8TO5(-28), .W8TO6(26), .W8TO7(-21), .W8TO8(324), .W8TO9(-82), .W9TO0(104), .W9TO1(-214), .W9TO2(162), .W9TO3(-151), .W9TO4(-252), .W9TO5(-155), .W9TO6(-117), .W9TO7(-185), .W9TO8(44), .W9TO9(176), .W10TO0(-74), .W10TO1(12), .W10TO2(117), .W10TO3(-72), .W10TO4(-173), .W10TO5(19), .W10TO6(79), .W10TO7(153), .W10TO8(-224), .W10TO9(-264), .W11TO0(-132), .W11TO1(110), .W11TO2(-77), .W11TO3(-80), .W11TO4(-210), .W11TO5(-10), .W11TO6(9), .W11TO7(-106), .W11TO8(-118), .W11TO9(87), .W12TO0(-114), .W12TO1(59), .W12TO2(-139), .W12TO3(156), .W12TO4(135), .W12TO5(-126), .W12TO6(-367), .W12TO7(165), .W12TO8(166), .W12TO9(-164), .W13TO0(87), .W13TO1(130), .W13TO2(193), .W13TO3(-87), .W13TO4(-299), .W13TO5(-260), .W13TO6(-161), .W13TO7(202), .W13TO8(129), .W13TO9(-139), .W14TO0(-110), .W14TO1(-137), .W14TO2(-3), .W14TO3(31), .W14TO4(62), .W14TO5(100), .W14TO6(-190), .W14TO7(94), .W14TO8(-179), .W14TO9(1), .W15TO0(22), .W15TO1(-247), .W15TO2(129), .W15TO3(36), .W15TO4(-126), .W15TO5(-273), .W15TO6(-100), .W15TO7(-88), .W15TO8(155), .W15TO9(195), .W16TO0(-18), .W16TO1(-159), .W16TO2(-265), .W16TO3(-245), .W16TO4(142), .W16TO5(174), .W16TO6(40), .W16TO7(72), .W16TO8(-78), .W16TO9(70), .W17TO0(-238), .W17TO1(361), .W17TO2(39), .W17TO3(1), .W17TO4(38), .W17TO5(-73), .W17TO6(-316), .W17TO7(204), .W17TO8(172), .W17TO9(-241), .W18TO0(-307), .W18TO1(-38), .W18TO2(15), .W18TO3(84), .W18TO4(-94), .W18TO5(243), .W18TO6(-26), .W18TO7(-174), .W18TO8(-137), .W18TO9(94), .W19TO0(-109), .W19TO1(-21), .W19TO2(299), .W19TO3(403), .W19TO4(-235), .W19TO5(-243), .W19TO6(-141), .W19TO7(-185), .W19TO8(54), .W19TO9(-37), .W20TO0(131), .W20TO1(-57), .W20TO2(-112), .W20TO3(-174), .W20TO4(179), .W20TO5(214), .W20TO6(-168), .W20TO7(66), .W20TO8(226), .W20TO9(-228), .W21TO0(-24), .W21TO1(55), .W21TO2(31), .W21TO3(-164), .W21TO4(-187), .W21TO5(75), .W21TO6(250), .W21TO7(128), .W21TO8(49), .W21TO9(-141), .W22TO0(82), .W22TO1(242), .W22TO2(154), .W22TO3(28), .W22TO4(-175), .W22TO5(-214), .W22TO6(112), .W22TO7(-223), .W22TO8(45), .W22TO9(205), .W23TO0(280), .W23TO1(-39), .W23TO2(77), .W23TO3(198), .W23TO4(-178), .W23TO5(224), .W23TO6(-44), .W23TO7(-50), .W23TO8(228), .W23TO9(59), .W24TO0(-152), .W24TO1(-197), .W24TO2(225), .W24TO3(78), .W24TO4(-246), .W24TO5(-149), .W24TO6(-157), .W24TO7(191), .W24TO8(153), .W24TO9(169), .W25TO0(-35), .W25TO1(229), .W25TO2(12), .W25TO3(149), .W25TO4(159), .W25TO5(76), .W25TO6(61), .W25TO7(-27), .W25TO8(-169), .W25TO9(-11), .W26TO0(199), .W26TO1(57), .W26TO2(-156), .W26TO3(174), .W26TO4(-108), .W26TO5(-30), .W26TO6(-18), .W26TO7(115), .W26TO8(-34), .W26TO9(219), .W27TO0(226), .W27TO1(8), .W27TO2(-30), .W27TO3(65), .W27TO4(13), .W27TO5(-66), .W27TO6(39), .W27TO7(147), .W27TO8(274), .W27TO9(230), .W28TO0(-120), .W28TO1(-53), .W28TO2(78), .W28TO3(60), .W28TO4(-169), .W28TO5(-95), .W28TO6(-73), .W28TO7(227), .W28TO8(161), .W28TO9(165), .W29TO0(266), .W29TO1(-447), .W29TO2(-7), .W29TO3(-133), .W29TO4(361), .W29TO5(-72), .W29TO6(-176), .W29TO7(321), .W29TO8(38), .W29TO9(291), .W30TO0(135), .W30TO1(-119), .W30TO2(-91), .W30TO3(-72), .W30TO4(-18), .W30TO5(-210), .W30TO6(344), .W30TO7(-63), .W30TO8(254), .W30TO9(15), .W31TO0(-150), .W31TO1(-54), .W31TO2(-129), .W31TO3(-103), .W31TO4(286), .W31TO5(-157), .W31TO6(114), .W31TO7(-30), .W31TO8(181), .W31TO9(-297), .W32TO0(-25), .W32TO1(-160), .W32TO2(-183), .W32TO3(-130), .W32TO4(160), .W32TO5(-236), .W32TO6(126), .W32TO7(-112), .W32TO8(-291), .W32TO9(-156), .W33TO0(92), .W33TO1(-195), .W33TO2(-286), .W33TO3(142), .W33TO4(96), .W33TO5(264), .W33TO6(230), .W33TO7(126), .W33TO8(202), .W33TO9(-187), .W34TO0(-89), .W34TO1(68), .W34TO2(-135), .W34TO3(-65), .W34TO4(-8), .W34TO5(214), .W34TO6(51), .W34TO7(-131), .W34TO8(63), .W34TO9(181), .W35TO0(87), .W35TO1(11), .W35TO2(-130), .W35TO3(-200), .W35TO4(-210), .W35TO5(41), .W35TO6(-3), .W35TO7(-190), .W35TO8(0), .W35TO9(178), .W36TO0(0), .W36TO1(55), .W36TO2(109), .W36TO3(-373), .W36TO4(136), .W36TO5(269), .W36TO6(116), .W36TO7(-214), .W36TO8(158), .W36TO9(-136), .W37TO0(-88), .W37TO1(137), .W37TO2(-91), .W37TO3(-81), .W37TO4(-260), .W37TO5(121), .W37TO6(-213), .W37TO7(-217), .W37TO8(-126), .W37TO9(12), .W38TO0(-40), .W38TO1(-169), .W38TO2(-107), .W38TO3(30), .W38TO4(40), .W38TO5(-228), .W38TO6(77), .W38TO7(-27), .W38TO8(-208), .W38TO9(-247), .W39TO0(-70), .W39TO1(-153), .W39TO2(37), .W39TO3(162), .W39TO4(288), .W39TO5(-166), .W39TO6(-14), .W39TO7(31), .W39TO8(-152), .W39TO9(136), .W40TO0(-168), .W40TO1(96), .W40TO2(242), .W40TO3(244), .W40TO4(69), .W40TO5(158), .W40TO6(238), .W40TO7(-92), .W40TO8(260), .W40TO9(160), .W41TO0(373), .W41TO1(-306), .W41TO2(139), .W41TO3(-87), .W41TO4(-111), .W41TO5(-211), .W41TO6(72), .W41TO7(-218), .W41TO8(249), .W41TO9(-256), .W42TO0(100), .W42TO1(231), .W42TO2(31), .W42TO3(223), .W42TO4(13), .W42TO5(170), .W42TO6(-123), .W42TO7(264), .W42TO8(215), .W42TO9(183), .W43TO0(-7), .W43TO1(167), .W43TO2(72), .W43TO3(131), .W43TO4(32), .W43TO5(-113), .W43TO6(-123), .W43TO7(-304), .W43TO8(50), .W43TO9(-52), .W44TO0(182), .W44TO1(-90), .W44TO2(112), .W44TO3(69), .W44TO4(-78), .W44TO5(-223), .W44TO6(-153), .W44TO7(-60), .W44TO8(-192), .W44TO9(165), .W45TO0(262), .W45TO1(101), .W45TO2(-135), .W45TO3(-30), .W45TO4(-176), .W45TO5(117), .W45TO6(219), .W45TO7(244), .W45TO8(119), .W45TO9(-50), .W46TO0(97), .W46TO1(0), .W46TO2(-34), .W46TO3(279), .W46TO4(198), .W46TO5(226), .W46TO6(-10), .W46TO7(83), .W46TO8(29), .W46TO9(235), .W47TO0(-211), .W47TO1(46), .W47TO2(55), .W47TO3(206), .W47TO4(-242), .W47TO5(-216), .W47TO6(-253), .W47TO7(189), .W47TO8(236), .W47TO9(359), .W48TO0(151), .W48TO1(-132), .W48TO2(29), .W48TO3(203), .W48TO4(76), .W48TO5(-180), .W48TO6(216), .W48TO7(-12), .W48TO8(-11), .W48TO9(191), .W49TO0(67), .W49TO1(27), .W49TO2(-446), .W49TO3(187), .W49TO4(-143), .W49TO5(15), .W49TO6(-89), .W49TO7(-292), .W49TO8(199), .W49TO9(-111), .W50TO0(-185), .W50TO1(-125), .W50TO2(107), .W50TO3(57), .W50TO4(43), .W50TO5(-163), .W50TO6(-72), .W50TO7(-99), .W50TO8(96), .W50TO9(135), .W51TO0(68), .W51TO1(-292), .W51TO2(-192), .W51TO3(-69), .W51TO4(150), .W51TO5(-202), .W51TO6(-47), .W51TO7(159), .W51TO8(105), .W51TO9(84), .W52TO0(-87), .W52TO1(-329), .W52TO2(164), .W52TO3(-130), .W52TO4(-246), .W52TO5(202), .W52TO6(131), .W52TO7(-82), .W52TO8(95), .W52TO9(-18), .W53TO0(-396), .W53TO1(129), .W53TO2(168), .W53TO3(-81), .W53TO4(-305), .W53TO5(96), .W53TO6(185), .W53TO7(54), .W53TO8(231), .W53TO9(-219), .W54TO0(44), .W54TO1(-230), .W54TO2(-253), .W54TO3(-221), .W54TO4(31), .W54TO5(42), .W54TO6(428), .W54TO7(94), .W54TO8(-71), .W54TO9(56), .W55TO0(-208), .W55TO1(220), .W55TO2(2), .W55TO3(-48), .W55TO4(-57), .W55TO5(-235), .W55TO6(129), .W55TO7(115), .W55TO8(4), .W55TO9(75), .W56TO0(-14), .W56TO1(-132), .W56TO2(-192), .W56TO3(-93), .W56TO4(-170), .W56TO5(138), .W56TO6(-106), .W56TO7(161), .W56TO8(-164), .W56TO9(-74), .W57TO0(225), .W57TO1(175), .W57TO2(166), .W57TO3(-170), .W57TO4(249), .W57TO5(-147), .W57TO6(50), .W57TO7(-41), .W57TO8(62), .W57TO9(-9), .W58TO0(192), .W58TO1(-49), .W58TO2(351), .W58TO3(-141), .W58TO4(86), .W58TO5(-44), .W58TO6(-2), .W58TO7(150), .W58TO8(181), .W58TO9(153), .W59TO0(314), .W59TO1(-218), .W59TO2(170), .W59TO3(51), .W59TO4(-97), .W59TO5(-73), .W59TO6(240), .W59TO7(53), .W59TO8(-320), .W59TO9(-392), .W60TO0(-212), .W60TO1(495), .W60TO2(-160), .W60TO3(-267), .W60TO4(266), .W60TO5(-120), .W60TO6(199), .W60TO7(-104), .W60TO8(-248), .W60TO9(7), .W61TO0(76), .W61TO1(117), .W61TO2(-91), .W61TO3(75), .W61TO4(-162), .W61TO5(-299), .W61TO6(-74), .W61TO7(396), .W61TO8(220), .W61TO9(116), .W62TO0(-119), .W62TO1(-181), .W62TO2(64), .W62TO3(-44), .W62TO4(57), .W62TO5(84), .W62TO6(-120), .W62TO7(241), .W62TO8(278), .W62TO9(218), .W63TO0(220), .W63TO1(-241), .W63TO2(77), .W63TO3(4), .W63TO4(-352), .W63TO5(19), .W63TO6(-41), .W63TO7(-135), .W63TO8(-157), .W63TO9(-75), .W64TO0(-17), .W64TO1(-46), .W64TO2(320), .W64TO3(-170), .W64TO4(-64), .W64TO5(145), .W64TO6(-118), .W64TO7(-19), .W64TO8(-42), .W64TO9(-58), .W65TO0(-198), .W65TO1(208), .W65TO2(130), .W65TO3(-39), .W65TO4(289), .W65TO5(51), .W65TO6(-171), .W65TO7(-204), .W65TO8(-166), .W65TO9(-119), .W66TO0(260), .W66TO1(160), .W66TO2(209), .W66TO3(258), .W66TO4(179), .W66TO5(239), .W66TO6(7), .W66TO7(27), .W66TO8(-90), .W66TO9(-30), .W67TO0(-139), .W67TO1(-101), .W67TO2(336), .W67TO3(232), .W67TO4(-76), .W67TO5(44), .W67TO6(144), .W67TO7(-102), .W67TO8(-323), .W67TO9(-224), .W68TO0(-121), .W68TO1(-102), .W68TO2(-264), .W68TO3(-209), .W68TO4(-179), .W68TO5(69), .W68TO6(58), .W68TO7(-243), .W68TO8(-270), .W68TO9(-206), .W69TO0(-22), .W69TO1(-125), .W69TO2(156), .W69TO3(140), .W69TO4(103), .W69TO5(70), .W69TO6(-207), .W69TO7(162), .W69TO8(-201), .W69TO9(-125), .W70TO0(-121), .W70TO1(-157), .W70TO2(154), .W70TO3(-95), .W70TO4(-67), .W70TO5(-270), .W70TO6(272), .W70TO7(-181), .W70TO8(228), .W70TO9(274), .W71TO0(207), .W71TO1(-76), .W71TO2(-216), .W71TO3(223), .W71TO4(43), .W71TO5(-51), .W71TO6(-62), .W71TO7(13), .W71TO8(26), .W71TO9(193), .W72TO0(163), .W72TO1(-88), .W72TO2(-202), .W72TO3(-131), .W72TO4(-116), .W72TO5(-112), .W72TO6(-163), .W72TO7(-276), .W72TO8(-227), .W72TO9(33), .W73TO0(-172), .W73TO1(120), .W73TO2(219), .W73TO3(-116), .W73TO4(-128), .W73TO5(163), .W73TO6(-26), .W73TO7(66), .W73TO8(56), .W73TO9(-136), .W74TO0(-77), .W74TO1(-16), .W74TO2(205), .W74TO3(224), .W74TO4(260), .W74TO5(186), .W74TO6(0), .W74TO7(223), .W74TO8(-65), .W74TO9(-13), .W75TO0(76), .W75TO1(54), .W75TO2(-186), .W75TO3(89), .W75TO4(6), .W75TO5(221), .W75TO6(137), .W75TO7(-135), .W75TO8(182), .W75TO9(182), .W76TO0(100), .W76TO1(-72), .W76TO2(120), .W76TO3(201), .W76TO4(-54), .W76TO5(112), .W76TO6(-35), .W76TO7(-256), .W76TO8(-67), .W76TO9(-266), .W77TO0(-9), .W77TO1(23), .W77TO2(-78), .W77TO3(-21), .W77TO4(-20), .W77TO5(244), .W77TO6(-14), .W77TO7(177), .W77TO8(104), .W77TO9(0), .W78TO0(21), .W78TO1(128), .W78TO2(206), .W78TO3(-295), .W78TO4(170), .W78TO5(-227), .W78TO6(-44), .W78TO7(195), .W78TO8(-341), .W78TO9(-401), .W79TO0(169), .W79TO1(6), .W79TO2(-60), .W79TO3(291), .W79TO4(-22), .W79TO5(61), .W79TO6(13), .W79TO7(26), .W79TO8(-111), .W79TO9(-256), .W80TO0(200), .W80TO1(56), .W80TO2(143), .W80TO3(-125), .W80TO4(84), .W80TO5(-231), .W80TO6(80), .W80TO7(-208), .W80TO8(396), .W80TO9(-165), .W81TO0(30), .W81TO1(-185), .W81TO2(-150), .W81TO3(-115), .W81TO4(-257), .W81TO5(3), .W81TO6(-72), .W81TO7(-131), .W81TO8(24), .W81TO9(-216), .W82TO0(-353), .W82TO1(97), .W82TO2(78), .W82TO3(165), .W82TO4(-320), .W82TO5(183), .W82TO6(260), .W82TO7(-358), .W82TO8(249), .W82TO9(292), .W83TO0(-29), .W83TO1(-234), .W83TO2(38), .W83TO3(362), .W83TO4(-83), .W83TO5(167), .W83TO6(-264), .W83TO7(-46), .W83TO8(-259), .W83TO9(320), .W84TO0(-177), .W84TO1(354), .W84TO2(-40), .W84TO3(-360), .W84TO4(217), .W84TO5(-267), .W84TO6(52), .W84TO7(88), .W84TO8(144), .W84TO9(250), .W85TO0(-174), .W85TO1(127), .W85TO2(-205), .W85TO3(-72), .W85TO4(-131), .W85TO5(-227), .W85TO6(-11), .W85TO7(112), .W85TO8(-225), .W85TO9(80), .W86TO0(27), .W86TO1(234), .W86TO2(-152), .W86TO3(132), .W86TO4(80), .W86TO5(6), .W86TO6(-150), .W86TO7(-51), .W86TO8(-231), .W86TO9(199), .W87TO0(248), .W87TO1(-222), .W87TO2(-136), .W87TO3(-153), .W87TO4(149), .W87TO5(225), .W87TO6(25), .W87TO7(-63), .W87TO8(171), .W87TO9(-41), .W88TO0(-153), .W88TO1(347), .W88TO2(-233), .W88TO3(39), .W88TO4(-13), .W88TO5(-162), .W88TO6(195), .W88TO7(3), .W88TO8(76), .W88TO9(135), .W89TO0(72), .W89TO1(250), .W89TO2(159), .W89TO3(-119), .W89TO4(-408), .W89TO5(-128), .W89TO6(163), .W89TO7(-142), .W89TO8(77), .W89TO9(-184), .W90TO0(-96), .W90TO1(159), .W90TO2(-49), .W90TO3(-217), .W90TO4(-61), .W90TO5(-170), .W90TO6(-247), .W90TO7(-212), .W90TO8(-117), .W90TO9(-226), .W91TO0(154), .W91TO1(80), .W91TO2(-26), .W91TO3(400), .W91TO4(-37), .W91TO5(-227), .W91TO6(-32), .W91TO7(-151), .W91TO8(-44), .W91TO9(-124), .W92TO0(-142), .W92TO1(84), .W92TO2(115), .W92TO3(6), .W92TO4(91), .W92TO5(46), .W92TO6(54), .W92TO7(149), .W92TO8(120), .W92TO9(-3), .W93TO0(-319), .W93TO1(20), .W93TO2(60), .W93TO3(176), .W93TO4(191), .W93TO5(-123), .W93TO6(144), .W93TO7(244), .W93TO8(213), .W93TO9(-378), .W94TO0(20), .W94TO1(152), .W94TO2(210), .W94TO3(129), .W94TO4(187), .W94TO5(-165), .W94TO6(235), .W94TO7(252), .W94TO8(23), .W94TO9(102), .W95TO0(-219), .W95TO1(83), .W95TO2(93), .W95TO3(245), .W95TO4(123), .W95TO5(-241), .W95TO6(79), .W95TO7(20), .W95TO8(2), .W95TO9(-338), .W96TO0(-119), .W96TO1(-29), .W96TO2(162), .W96TO3(-34), .W96TO4(-13), .W96TO5(48), .W96TO6(-233), .W96TO7(33), .W96TO8(141), .W96TO9(-121), .W97TO0(231), .W97TO1(-51), .W97TO2(1), .W97TO3(-19), .W97TO4(-174), .W97TO5(-38), .W97TO6(-29), .W97TO7(65), .W97TO8(-79), .W97TO9(-106), .W98TO0(-26), .W98TO1(7), .W98TO2(155), .W98TO3(-145), .W98TO4(147), .W98TO5(-264), .W98TO6(24), .W98TO7(-342), .W98TO8(91), .W98TO9(89), .W99TO0(-179), .W99TO1(-280), .W99TO2(-261), .W99TO3(-132), .W99TO4(85), .W99TO5(1), .W99TO6(-65), .W99TO7(1), .W99TO8(140), .W99TO9(-196)) layer1(.clk(clk), .rst(rst), .in0(con0[0]), .in1(con0[1]), .in2(con0[2]), .in3(con0[3]), .in4(con0[4]), .in5(con0[5]), .in6(con0[6]), .in7(con0[7]), .in8(con0[8]), .in9(con0[9]), .in10(con0[10]), .in11(con0[11]), .in12(con0[12]), .in13(con0[13]), .in14(con0[14]), .in15(con0[15]), .in16(con0[16]), .in17(con0[17]), .in18(con0[18]), .in19(con0[19]), .in20(con0[20]), .in21(con0[21]), .in22(con0[22]), .in23(con0[23]), .in24(con0[24]), .in25(con0[25]), .in26(con0[26]), .in27(con0[27]), .in28(con0[28]), .in29(con0[29]), .in30(con0[30]), .in31(con0[31]), .in32(con0[32]), .in33(con0[33]), .in34(con0[34]), .in35(con0[35]), .in36(con0[36]), .in37(con0[37]), .in38(con0[38]), .in39(con0[39]), .in40(con0[40]), .in41(con0[41]), .in42(con0[42]), .in43(con0[43]), .in44(con0[44]), .in45(con0[45]), .in46(con0[46]), .in47(con0[47]), .in48(con0[48]), .in49(con0[49]), .in50(con0[50]), .in51(con0[51]), .in52(con0[52]), .in53(con0[53]), .in54(con0[54]), .in55(con0[55]), .in56(con0[56]), .in57(con0[57]), .in58(con0[58]), .in59(con0[59]), .in60(con0[60]), .in61(con0[61]), .in62(con0[62]), .in63(con0[63]), .in64(con0[64]), .in65(con0[65]), .in66(con0[66]), .in67(con0[67]), .in68(con0[68]), .in69(con0[69]), .in70(con0[70]), .in71(con0[71]), .in72(con0[72]), .in73(con0[73]), .in74(con0[74]), .in75(con0[75]), .in76(con0[76]), .in77(con0[77]), .in78(con0[78]), .in79(con0[79]), .in80(con0[80]), .in81(con0[81]), .in82(con0[82]), .in83(con0[83]), .in84(con0[84]), .in85(con0[85]), .in86(con0[86]), .in87(con0[87]), .in88(con0[88]), .in89(con0[89]), .in90(con0[90]), .in91(con0[91]), .in92(con0[92]), .in93(con0[93]), .in94(con0[94]), .in95(con0[95]), .in96(con0[96]), .in97(con0[97]), .in98(con0[98]), .in99(con0[99]), .out0(out0), .out1(out1), .out2(out2), .out3(out3), .out4(out4), .out5(out5), .out6(out6), .out7(out7), .out8(out8), .out9(out9));

endmodule

module testbench_digits;

logic clk;
logic rst;

reg [15:0] net_in0, net_in1, net_in2, net_in3, net_in4, net_in5, net_in6, net_in7, net_in8, net_in9, net_in10, net_in11, net_in12, net_in13, net_in14, net_in15, net_in16, net_in17, net_in18, net_in19, net_in20, net_in21, net_in22, net_in23, net_in24, net_in25, net_in26, net_in27, net_in28, net_in29, net_in30, net_in31, net_in32, net_in33, net_in34, net_in35, net_in36, net_in37, net_in38, net_in39, net_in40, net_in41, net_in42, net_in43, net_in44, net_in45, net_in46, net_in47, net_in48, net_in49, net_in50, net_in51, net_in52, net_in53, net_in54, net_in55, net_in56, net_in57, net_in58, net_in59, net_in60, net_in61, net_in62, net_in63;
wire [15:0] net_out0, net_out1, net_out2, net_out3, net_out4, net_out5, net_out6, net_out7, net_out8, net_out9;

network net(.clk(clk), .rst(rst), .in0(net_in0), .in1(net_in1), .in2(net_in2), .in3(net_in3), .in4(net_in4), .in5(net_in5), .in6(net_in6), .in7(net_in7), .in8(net_in8), .in9(net_in9), .in10(net_in10), .in11(net_in11), .in12(net_in12), .in13(net_in13), .in14(net_in14), .in15(net_in15), .in16(net_in16), .in17(net_in17), .in18(net_in18), .in19(net_in19), .in20(net_in20), .in21(net_in21), .in22(net_in22), .in23(net_in23), .in24(net_in24), .in25(net_in25), .in26(net_in26), .in27(net_in27), .in28(net_in28), .in29(net_in29), .in30(net_in30), .in31(net_in31), .in32(net_in32), .in33(net_in33), .in34(net_in34), .in35(net_in35), .in36(net_in36), .in37(net_in37), .in38(net_in38), .in39(net_in39), .in40(net_in40), .in41(net_in41), .in42(net_in42), .in43(net_in43), .in44(net_in44), .in45(net_in45), .in46(net_in46), .in47(net_in47), .in48(net_in48), .in49(net_in49), .in50(net_in50), .in51(net_in51), .in52(net_in52), .in53(net_in53), .in54(net_in54), .in55(net_in55), .in56(net_in56), .in57(net_in57), .in58(net_in58), .in59(net_in59), .in60(net_in60), .in61(net_in61), .in62(net_in62), .in63(net_in63), .out0(net_out0), .out1(net_out1), .out2(net_out2), .out3(net_out3), .out4(net_out4), .out5(net_out5), .out6(net_out6), .out7(net_out7), .out8(net_out8), .out9(net_out9));

task test;
input [15:0] in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63;
begin
    net_in0 = in0;
    net_in1 = in1;
    net_in2 = in2;
    net_in3 = in3;
    net_in4 = in4;
    net_in5 = in5;
    net_in6 = in6;
    net_in7 = in7;
    net_in8 = in8;
    net_in9 = in9;
    net_in10 = in10;
    net_in11 = in11;
    net_in12 = in12;
    net_in13 = in13;
    net_in14 = in14;
    net_in15 = in15;
    net_in16 = in16;
    net_in17 = in17;
    net_in18 = in18;
    net_in19 = in19;
    net_in20 = in20;
    net_in21 = in21;
    net_in22 = in22;
    net_in23 = in23;
    net_in24 = in24;
    net_in25 = in25;
    net_in26 = in26;
    net_in27 = in27;
    net_in28 = in28;
    net_in29 = in29;
    net_in30 = in30;
    net_in31 = in31;
    net_in32 = in32;
    net_in33 = in33;
    net_in34 = in34;
    net_in35 = in35;
    net_in36 = in36;
    net_in37 = in37;
    net_in38 = in38;
    net_in39 = in39;
    net_in40 = in40;
    net_in41 = in41;
    net_in42 = in42;
    net_in43 = in43;
    net_in44 = in44;
    net_in45 = in45;
    net_in46 = in46;
    net_in47 = in47;
    net_in48 = in48;
    net_in49 = in49;
    net_in50 = in50;
    net_in51 = in51;
    net_in52 = in52;
    net_in53 = in53;
    net_in54 = in54;
    net_in55 = in55;
    net_in56 = in56;
    net_in57 = in57;
    net_in58 = in58;
    net_in59 = in59;
    net_in60 = in60;
    net_in61 = in61;
    net_in62 = in62;
    net_in63 = in63;
    #10000000

    $write("%d ", net_out0);
    $write("%d ", net_out1);
    $write("%d ", net_out2);
    $write("%d ", net_out3);
    $write("%d ", net_out4);
    $write("%d ", net_out5);
    $write("%d ", net_out6);
    $write("%d ", net_out7);
    $write("%d ", net_out8);
    $write("%d ", net_out9);
    $display();
end
endtask

initial begin
    test(0, 0, 1000, 15000, 15000, 2000, 0, 0, 0, 0, 3000, 12000, 16000, 6000, 0, 0, 0, 0, 0, 4000, 16000, 4000, 0, 0, 0, 0, 3000, 8000, 16000, 4000, 0, 0, 0, 10000, 16000, 16000, 16000, 16000, 8000, 0, 0, 8000, 11000, 14000, 14000, 5000, 1000, 0, 0, 0, 0, 15000, 6000, 0, 0, 0, 0, 0, 1000, 15000, 2000, 0, 0, 0);
    test(0, 0, 13000, 13000, 8000, 2000, 0, 0, 0, 5000, 16000, 16000, 16000, 12000, 0, 0, 0, 1000, 15000, 12000, 0, 0, 0, 0, 0, 0, 12000, 13000, 7000, 1000, 0, 0, 0, 0, 8000, 16000, 16000, 12000, 0, 0, 0, 0, 0, 4000, 9000, 16000, 3000, 0, 0, 0, 1000, 5000, 14000, 15000, 1000, 0, 0, 0, 10000, 16000, 16000, 6000, 0, 0);
    test(0, 0, 14000, 12000, 12000, 12000, 6000, 0, 0, 2000, 15000, 8000, 8000, 8000, 4000, 0, 0, 5000, 12000, 0, 0, 0, 0, 0, 0, 8000, 16000, 12000, 11000, 7000, 0, 0, 0, 1000, 4000, 4000, 9000, 15000, 7000, 0, 0, 0, 0, 0, 0, 8000, 8000, 0, 0, 1000, 11000, 4000, 5000, 14000, 7000, 0, 0, 0, 12000, 16000, 16000, 8000, 1000, 0);
    test(0, 0, 0, 5000, 13000, 16000, 8000, 0, 0, 0, 8000, 15000, 6000, 7000, 14000, 0, 0, 2000, 16000, 1000, 1000, 11000, 10000, 0, 0, 4000, 16000, 15000, 16000, 16000, 6000, 0, 0, 0, 4000, 4000, 5000, 15000, 1000, 0, 0, 0, 0, 0, 9000, 8000, 0, 0, 0, 0, 0, 2000, 15000, 1000, 0, 0, 0, 0, 0, 6000, 10000, 0, 0, 0);
    test(0, 0, 5000, 13000, 16000, 14000, 0, 0, 0, 1000, 14000, 8000, 5000, 16000, 2000, 0, 0, 0, 1000, 0, 2000, 15000, 2000, 0, 0, 0, 0, 2000, 8000, 15000, 3000, 0, 0, 0, 0, 15000, 16000, 13000, 8000, 0, 0, 0, 0, 6000, 14000, 0, 0, 0, 0, 0, 0, 13000, 7000, 0, 0, 0, 0, 0, 7000, 14000, 0, 0, 0, 0);
    test(0, 2000, 13000, 16000, 16000, 16000, 15000, 2000, 0, 8000, 16000, 12000, 8000, 4000, 1000, 0, 0, 5000, 16000, 13000, 1000, 0, 0, 0, 0, 0, 8000, 16000, 8000, 0, 0, 0, 0, 0, 0, 10000, 16000, 0, 0, 0, 0, 0, 0, 9000, 16000, 0, 0, 0, 0, 0, 3000, 13000, 12000, 0, 0, 0, 0, 2000, 16000, 16000, 6000, 0, 0, 0);
    test(0, 1000, 12000, 15000, 16000, 13000, 1000, 0, 0, 4000, 16000, 15000, 7000, 15000, 4000, 0, 0, 0, 16000, 6000, 11000, 15000, 2000, 0, 0, 0, 9000, 16000, 15000, 4000, 0, 0, 0, 0, 8000, 16000, 8000, 0, 0, 0, 0, 0, 15000, 15000, 11000, 0, 0, 0, 0, 2000, 16000, 10000, 12000, 0, 0, 0, 0, 2000, 13000, 16000, 10000, 0, 0, 0);
    test(0, 3000, 12000, 12000, 14000, 4000, 0, 0, 0, 1000, 13000, 4000, 4000, 0, 0, 0, 0, 4000, 14000, 4000, 3000, 0, 0, 0, 0, 5000, 13000, 12000, 14000, 10000, 0, 0, 0, 0, 0, 0, 0, 11000, 6000, 0, 0, 0, 0, 0, 0, 4000, 8000, 0, 0, 0, 6000, 2000, 0, 8000, 8000, 0, 0, 2000, 13000, 16000, 16000, 16000, 2000, 0);
    test(0, 0, 4000, 14000, 16000, 5000, 0, 0, 0, 4000, 16000, 16000, 16000, 8000, 0, 0, 0, 12000, 12000, 0, 15000, 8000, 0, 0, 0, 2000, 1000, 5000, 16000, 13000, 1000, 0, 0, 0, 0, 1000, 11000, 15000, 11000, 0, 0, 0, 0, 0, 0, 11000, 12000, 0, 0, 0, 2000, 13000, 12000, 16000, 7000, 0, 0, 0, 3000, 16000, 15000, 8000, 0, 0);
    test(0, 0, 5000, 8000, 11000, 5000, 0, 0, 0, 0, 13000, 16000, 12000, 12000, 0, 0, 0, 1000, 16000, 9000, 0, 9000, 3000, 0, 0, 3000, 16000, 6000, 0, 6000, 6000, 0, 0, 3000, 11000, 1000, 0, 5000, 6000, 0, 0, 0, 12000, 0, 0, 11000, 6000, 0, 0, 0, 14000, 5000, 12000, 15000, 1000, 0, 0, 0, 6000, 16000, 13000, 2000, 0, 0);
end
endmodule
