module neuron65in(clk, rst, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, out);

parameter signed BIAS = 0;
parameter signed W0 = 0;
parameter signed W1 = 0;
parameter signed W2 = 0;
parameter signed W3 = 0;
parameter signed W4 = 0;
parameter signed W5 = 0;
parameter signed W6 = 0;
parameter signed W7 = 0;
parameter signed W8 = 0;
parameter signed W9 = 0;
parameter signed W10 = 0;
parameter signed W11 = 0;
parameter signed W12 = 0;
parameter signed W13 = 0;
parameter signed W14 = 0;
parameter signed W15 = 0;
parameter signed W16 = 0;
parameter signed W17 = 0;
parameter signed W18 = 0;
parameter signed W19 = 0;
parameter signed W20 = 0;
parameter signed W21 = 0;
parameter signed W22 = 0;
parameter signed W23 = 0;
parameter signed W24 = 0;
parameter signed W25 = 0;
parameter signed W26 = 0;
parameter signed W27 = 0;
parameter signed W28 = 0;
parameter signed W29 = 0;
parameter signed W30 = 0;
parameter signed W31 = 0;
parameter signed W32 = 0;
parameter signed W33 = 0;
parameter signed W34 = 0;
parameter signed W35 = 0;
parameter signed W36 = 0;
parameter signed W37 = 0;
parameter signed W38 = 0;
parameter signed W39 = 0;
parameter signed W40 = 0;
parameter signed W41 = 0;
parameter signed W42 = 0;
parameter signed W43 = 0;
parameter signed W44 = 0;
parameter signed W45 = 0;
parameter signed W46 = 0;
parameter signed W47 = 0;
parameter signed W48 = 0;
parameter signed W49 = 0;
parameter signed W50 = 0;
parameter signed W51 = 0;
parameter signed W52 = 0;
parameter signed W53 = 0;
parameter signed W54 = 0;
parameter signed W55 = 0;
parameter signed W56 = 0;
parameter signed W57 = 0;
parameter signed W58 = 0;
parameter signed W59 = 0;
parameter signed W60 = 0;
parameter signed W61 = 0;
parameter signed W62 = 0;
parameter signed W63 = 0;
parameter signed W64 = 0;

input wire clk;
input wire rst;

input signed [63:0] in0;
input signed [63:0] in1;
input signed [63:0] in2;
input signed [63:0] in3;
input signed [63:0] in4;
input signed [63:0] in5;
input signed [63:0] in6;
input signed [63:0] in7;
input signed [63:0] in8;
input signed [63:0] in9;
input signed [63:0] in10;
input signed [63:0] in11;
input signed [63:0] in12;
input signed [63:0] in13;
input signed [63:0] in14;
input signed [63:0] in15;
input signed [63:0] in16;
input signed [63:0] in17;
input signed [63:0] in18;
input signed [63:0] in19;
input signed [63:0] in20;
input signed [63:0] in21;
input signed [63:0] in22;
input signed [63:0] in23;
input signed [63:0] in24;
input signed [63:0] in25;
input signed [63:0] in26;
input signed [63:0] in27;
input signed [63:0] in28;
input signed [63:0] in29;
input signed [63:0] in30;
input signed [63:0] in31;
input signed [63:0] in32;
input signed [63:0] in33;
input signed [63:0] in34;
input signed [63:0] in35;
input signed [63:0] in36;
input signed [63:0] in37;
input signed [63:0] in38;
input signed [63:0] in39;
input signed [63:0] in40;
input signed [63:0] in41;
input signed [63:0] in42;
input signed [63:0] in43;
input signed [63:0] in44;
input signed [63:0] in45;
input signed [63:0] in46;
input signed [63:0] in47;
input signed [63:0] in48;
input signed [63:0] in49;
input signed [63:0] in50;
input signed [63:0] in51;
input signed [63:0] in52;
input signed [63:0] in53;
input signed [63:0] in54;
input signed [63:0] in55;
input signed [63:0] in56;
input signed [63:0] in57;
input signed [63:0] in58;
input signed [63:0] in59;
input signed [63:0] in60;
input signed [63:0] in61;
input signed [63:0] in62;
input signed [63:0] in63;
input signed [63:0] in64;

output reg signed [63:0] out;

reg signed [191:0] x;
reg signed [191:0] abs_x;
reg signed [191:0] y;
reg signed [191:0] sum_0_0;
reg signed [191:0] sum_0_1;
reg signed [191:0] sum_0_2;
reg signed [191:0] sum_0_3;
reg signed [191:0] sum_0_4;
reg signed [191:0] sum_0_5;
reg signed [191:0] sum_0_6;
reg signed [191:0] sum_0_7;
reg signed [191:0] sum_0_8;
reg signed [191:0] sum_0_9;
reg signed [191:0] sum_0_10;
reg signed [191:0] sum_0_11;
reg signed [191:0] sum_0_12;
reg signed [191:0] sum_0_13;
reg signed [191:0] sum_0_14;
reg signed [191:0] sum_0_15;
reg signed [191:0] sum_0_16;
reg signed [191:0] sum_0_17;
reg signed [191:0] sum_0_18;
reg signed [191:0] sum_0_19;
reg signed [191:0] sum_0_20;
reg signed [191:0] sum_0_21;
reg signed [191:0] sum_0_22;
reg signed [191:0] sum_0_23;
reg signed [191:0] sum_0_24;
reg signed [191:0] sum_0_25;
reg signed [191:0] sum_0_26;
reg signed [191:0] sum_0_27;
reg signed [191:0] sum_0_28;
reg signed [191:0] sum_0_29;
reg signed [191:0] sum_0_30;
reg signed [191:0] sum_0_31;
reg signed [191:0] sum_0_32;
reg signed [191:0] sum_1_0;
reg signed [191:0] sum_1_1;
reg signed [191:0] sum_1_2;
reg signed [191:0] sum_1_3;
reg signed [191:0] sum_1_4;
reg signed [191:0] sum_1_5;
reg signed [191:0] sum_1_6;
reg signed [191:0] sum_1_7;
reg signed [191:0] sum_1_8;
reg signed [191:0] sum_1_9;
reg signed [191:0] sum_1_10;
reg signed [191:0] sum_1_11;
reg signed [191:0] sum_1_12;
reg signed [191:0] sum_1_13;
reg signed [191:0] sum_1_14;
reg signed [191:0] sum_1_15;
reg signed [191:0] sum_2_0;
reg signed [191:0] sum_2_1;
reg signed [191:0] sum_2_2;
reg signed [191:0] sum_2_3;
reg signed [191:0] sum_2_4;
reg signed [191:0] sum_2_5;
reg signed [191:0] sum_2_6;
reg signed [191:0] sum_2_7;
reg signed [191:0] sum_3_0;
reg signed [191:0] sum_3_1;
reg signed [191:0] sum_3_2;
reg signed [191:0] sum_3_3;
reg signed [191:0] sum_4_0;
reg signed [191:0] sum_4_1;
reg signed [191:0] sum_5_0;
always @* begin
    sum_0_0 <= (in0 * W0 + 500000) / 1000000 + (in1 * W1 + 500000) / 1000000;
    sum_0_1 <= (in2 * W2 + 500000) / 1000000 + (in3 * W3 + 500000) / 1000000;
    sum_0_2 <= (in4 * W4 + 500000) / 1000000 + (in5 * W5 + 500000) / 1000000;
    sum_0_3 <= (in6 * W6 + 500000) / 1000000 + (in7 * W7 + 500000) / 1000000;
    sum_0_4 <= (in8 * W8 + 500000) / 1000000 + (in9 * W9 + 500000) / 1000000;
    sum_0_5 <= (in10 * W10 + 500000) / 1000000 + (in11 * W11 + 500000) / 1000000;
    sum_0_6 <= (in12 * W12 + 500000) / 1000000 + (in13 * W13 + 500000) / 1000000;
    sum_0_7 <= (in14 * W14 + 500000) / 1000000 + (in15 * W15 + 500000) / 1000000;
    sum_0_8 <= (in16 * W16 + 500000) / 1000000 + (in17 * W17 + 500000) / 1000000;
    sum_0_9 <= (in18 * W18 + 500000) / 1000000 + (in19 * W19 + 500000) / 1000000;
    sum_0_10 <= (in20 * W20 + 500000) / 1000000 + (in21 * W21 + 500000) / 1000000;
    sum_0_11 <= (in22 * W22 + 500000) / 1000000 + (in23 * W23 + 500000) / 1000000;
    sum_0_12 <= (in24 * W24 + 500000) / 1000000 + (in25 * W25 + 500000) / 1000000;
    sum_0_13 <= (in26 * W26 + 500000) / 1000000 + (in27 * W27 + 500000) / 1000000;
    sum_0_14 <= (in28 * W28 + 500000) / 1000000 + (in29 * W29 + 500000) / 1000000;
    sum_0_15 <= (in30 * W30 + 500000) / 1000000 + (in31 * W31 + 500000) / 1000000;
    sum_0_16 <= (in32 * W32 + 500000) / 1000000 + (in33 * W33 + 500000) / 1000000;
    sum_0_17 <= (in34 * W34 + 500000) / 1000000 + (in35 * W35 + 500000) / 1000000;
    sum_0_18 <= (in36 * W36 + 500000) / 1000000 + (in37 * W37 + 500000) / 1000000;
    sum_0_19 <= (in38 * W38 + 500000) / 1000000 + (in39 * W39 + 500000) / 1000000;
    sum_0_20 <= (in40 * W40 + 500000) / 1000000 + (in41 * W41 + 500000) / 1000000;
    sum_0_21 <= (in42 * W42 + 500000) / 1000000 + (in43 * W43 + 500000) / 1000000;
    sum_0_22 <= (in44 * W44 + 500000) / 1000000 + (in45 * W45 + 500000) / 1000000;
    sum_0_23 <= (in46 * W46 + 500000) / 1000000 + (in47 * W47 + 500000) / 1000000;
    sum_0_24 <= (in48 * W48 + 500000) / 1000000 + (in49 * W49 + 500000) / 1000000;
    sum_0_25 <= (in50 * W50 + 500000) / 1000000 + (in51 * W51 + 500000) / 1000000;
    sum_0_26 <= (in52 * W52 + 500000) / 1000000 + (in53 * W53 + 500000) / 1000000;
    sum_0_27 <= (in54 * W54 + 500000) / 1000000 + (in55 * W55 + 500000) / 1000000;
    sum_0_28 <= (in56 * W56 + 500000) / 1000000 + (in57 * W57 + 500000) / 1000000;
    sum_0_29 <= (in58 * W58 + 500000) / 1000000 + (in59 * W59 + 500000) / 1000000;
    sum_0_30 <= (in60 * W60 + 500000) / 1000000 + (in61 * W61 + 500000) / 1000000;
    sum_0_31 <= (in62 * W62 + 500000) / 1000000 + (in63 * W63 + 500000) / 1000000;
    sum_0_32 <= (in64 * W64 + 500000) / 1000000 + BIAS;
    sum_1_0 <= sum_0_0 + sum_0_1;
    sum_1_1 <= sum_0_2 + sum_0_3;
    sum_1_2 <= sum_0_4 + sum_0_5;
    sum_1_3 <= sum_0_6 + sum_0_7;
    sum_1_4 <= sum_0_8 + sum_0_9;
    sum_1_5 <= sum_0_10 + sum_0_11;
    sum_1_6 <= sum_0_12 + sum_0_13;
    sum_1_7 <= sum_0_14 + sum_0_15;
    sum_1_8 <= sum_0_16 + sum_0_17;
    sum_1_9 <= sum_0_18 + sum_0_19;
    sum_1_10 <= sum_0_20 + sum_0_21;
    sum_1_11 <= sum_0_22 + sum_0_23;
    sum_1_12 <= sum_0_24 + sum_0_25;
    sum_1_13 <= sum_0_26 + sum_0_27;
    sum_1_14 <= sum_0_28 + sum_0_29;
    sum_1_15 <= sum_0_30 + sum_0_31 + sum_0_32;
    sum_2_0 <= sum_1_0 + sum_1_1;
    sum_2_1 <= sum_1_2 + sum_1_3;
    sum_2_2 <= sum_1_4 + sum_1_5;
    sum_2_3 <= sum_1_6 + sum_1_7;
    sum_2_4 <= sum_1_8 + sum_1_9;
    sum_2_5 <= sum_1_10 + sum_1_11;
    sum_2_6 <= sum_1_12 + sum_1_13;
    sum_2_7 <= sum_1_14 + sum_1_15;
    sum_3_0 <= sum_2_0 + sum_2_1;
    sum_3_1 <= sum_2_2 + sum_2_3;
    sum_3_2 <= sum_2_4 + sum_2_5;
    sum_3_3 <= sum_2_6 + sum_2_7;
    sum_4_0 <= sum_3_0 + sum_3_1;
    sum_4_1 <= sum_3_2 + sum_3_3;
    sum_5_0 <= sum_4_0 + sum_4_1;
    x <= sum_5_0;
    abs_x = x < 0 ? -x : x;
    if (abs_x >= 5000000) y = 1000000;
    else if (abs_x >= 2375000) y = 31250 * abs_x / 1000000 + 843750;
    else if (abs_x >= 1000000) y = 125000 * abs_x / 1000000 + 625000;
    else y = 250000 * abs_x / 1000000 + 500000;
    out = x < 0 ? 1000000 - y : y;
end

endmodule

module neuron64in(clk, rst, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, out);

parameter signed BIAS = 0;
parameter signed W0 = 0;
parameter signed W1 = 0;
parameter signed W2 = 0;
parameter signed W3 = 0;
parameter signed W4 = 0;
parameter signed W5 = 0;
parameter signed W6 = 0;
parameter signed W7 = 0;
parameter signed W8 = 0;
parameter signed W9 = 0;
parameter signed W10 = 0;
parameter signed W11 = 0;
parameter signed W12 = 0;
parameter signed W13 = 0;
parameter signed W14 = 0;
parameter signed W15 = 0;
parameter signed W16 = 0;
parameter signed W17 = 0;
parameter signed W18 = 0;
parameter signed W19 = 0;
parameter signed W20 = 0;
parameter signed W21 = 0;
parameter signed W22 = 0;
parameter signed W23 = 0;
parameter signed W24 = 0;
parameter signed W25 = 0;
parameter signed W26 = 0;
parameter signed W27 = 0;
parameter signed W28 = 0;
parameter signed W29 = 0;
parameter signed W30 = 0;
parameter signed W31 = 0;
parameter signed W32 = 0;
parameter signed W33 = 0;
parameter signed W34 = 0;
parameter signed W35 = 0;
parameter signed W36 = 0;
parameter signed W37 = 0;
parameter signed W38 = 0;
parameter signed W39 = 0;
parameter signed W40 = 0;
parameter signed W41 = 0;
parameter signed W42 = 0;
parameter signed W43 = 0;
parameter signed W44 = 0;
parameter signed W45 = 0;
parameter signed W46 = 0;
parameter signed W47 = 0;
parameter signed W48 = 0;
parameter signed W49 = 0;
parameter signed W50 = 0;
parameter signed W51 = 0;
parameter signed W52 = 0;
parameter signed W53 = 0;
parameter signed W54 = 0;
parameter signed W55 = 0;
parameter signed W56 = 0;
parameter signed W57 = 0;
parameter signed W58 = 0;
parameter signed W59 = 0;
parameter signed W60 = 0;
parameter signed W61 = 0;
parameter signed W62 = 0;
parameter signed W63 = 0;

input wire clk;
input wire rst;

input signed [63:0] in0;
input signed [63:0] in1;
input signed [63:0] in2;
input signed [63:0] in3;
input signed [63:0] in4;
input signed [63:0] in5;
input signed [63:0] in6;
input signed [63:0] in7;
input signed [63:0] in8;
input signed [63:0] in9;
input signed [63:0] in10;
input signed [63:0] in11;
input signed [63:0] in12;
input signed [63:0] in13;
input signed [63:0] in14;
input signed [63:0] in15;
input signed [63:0] in16;
input signed [63:0] in17;
input signed [63:0] in18;
input signed [63:0] in19;
input signed [63:0] in20;
input signed [63:0] in21;
input signed [63:0] in22;
input signed [63:0] in23;
input signed [63:0] in24;
input signed [63:0] in25;
input signed [63:0] in26;
input signed [63:0] in27;
input signed [63:0] in28;
input signed [63:0] in29;
input signed [63:0] in30;
input signed [63:0] in31;
input signed [63:0] in32;
input signed [63:0] in33;
input signed [63:0] in34;
input signed [63:0] in35;
input signed [63:0] in36;
input signed [63:0] in37;
input signed [63:0] in38;
input signed [63:0] in39;
input signed [63:0] in40;
input signed [63:0] in41;
input signed [63:0] in42;
input signed [63:0] in43;
input signed [63:0] in44;
input signed [63:0] in45;
input signed [63:0] in46;
input signed [63:0] in47;
input signed [63:0] in48;
input signed [63:0] in49;
input signed [63:0] in50;
input signed [63:0] in51;
input signed [63:0] in52;
input signed [63:0] in53;
input signed [63:0] in54;
input signed [63:0] in55;
input signed [63:0] in56;
input signed [63:0] in57;
input signed [63:0] in58;
input signed [63:0] in59;
input signed [63:0] in60;
input signed [63:0] in61;
input signed [63:0] in62;
input signed [63:0] in63;

output reg signed [63:0] out;

reg signed [191:0] x;
reg signed [191:0] abs_x;
reg signed [191:0] y;
reg signed [191:0] sum_0_0;
reg signed [191:0] sum_0_1;
reg signed [191:0] sum_0_2;
reg signed [191:0] sum_0_3;
reg signed [191:0] sum_0_4;
reg signed [191:0] sum_0_5;
reg signed [191:0] sum_0_6;
reg signed [191:0] sum_0_7;
reg signed [191:0] sum_0_8;
reg signed [191:0] sum_0_9;
reg signed [191:0] sum_0_10;
reg signed [191:0] sum_0_11;
reg signed [191:0] sum_0_12;
reg signed [191:0] sum_0_13;
reg signed [191:0] sum_0_14;
reg signed [191:0] sum_0_15;
reg signed [191:0] sum_0_16;
reg signed [191:0] sum_0_17;
reg signed [191:0] sum_0_18;
reg signed [191:0] sum_0_19;
reg signed [191:0] sum_0_20;
reg signed [191:0] sum_0_21;
reg signed [191:0] sum_0_22;
reg signed [191:0] sum_0_23;
reg signed [191:0] sum_0_24;
reg signed [191:0] sum_0_25;
reg signed [191:0] sum_0_26;
reg signed [191:0] sum_0_27;
reg signed [191:0] sum_0_28;
reg signed [191:0] sum_0_29;
reg signed [191:0] sum_0_30;
reg signed [191:0] sum_0_31;
reg signed [191:0] sum_1_0;
reg signed [191:0] sum_1_1;
reg signed [191:0] sum_1_2;
reg signed [191:0] sum_1_3;
reg signed [191:0] sum_1_4;
reg signed [191:0] sum_1_5;
reg signed [191:0] sum_1_6;
reg signed [191:0] sum_1_7;
reg signed [191:0] sum_1_8;
reg signed [191:0] sum_1_9;
reg signed [191:0] sum_1_10;
reg signed [191:0] sum_1_11;
reg signed [191:0] sum_1_12;
reg signed [191:0] sum_1_13;
reg signed [191:0] sum_1_14;
reg signed [191:0] sum_1_15;
reg signed [191:0] sum_2_0;
reg signed [191:0] sum_2_1;
reg signed [191:0] sum_2_2;
reg signed [191:0] sum_2_3;
reg signed [191:0] sum_2_4;
reg signed [191:0] sum_2_5;
reg signed [191:0] sum_2_6;
reg signed [191:0] sum_2_7;
reg signed [191:0] sum_3_0;
reg signed [191:0] sum_3_1;
reg signed [191:0] sum_3_2;
reg signed [191:0] sum_3_3;
reg signed [191:0] sum_4_0;
reg signed [191:0] sum_4_1;
reg signed [191:0] sum_5_0;
always @* begin
    sum_0_0 <= (in0 * W0 + 500000) / 1000000 + (in1 * W1 + 500000) / 1000000;
    sum_0_1 <= (in2 * W2 + 500000) / 1000000 + (in3 * W3 + 500000) / 1000000;
    sum_0_2 <= (in4 * W4 + 500000) / 1000000 + (in5 * W5 + 500000) / 1000000;
    sum_0_3 <= (in6 * W6 + 500000) / 1000000 + (in7 * W7 + 500000) / 1000000;
    sum_0_4 <= (in8 * W8 + 500000) / 1000000 + (in9 * W9 + 500000) / 1000000;
    sum_0_5 <= (in10 * W10 + 500000) / 1000000 + (in11 * W11 + 500000) / 1000000;
    sum_0_6 <= (in12 * W12 + 500000) / 1000000 + (in13 * W13 + 500000) / 1000000;
    sum_0_7 <= (in14 * W14 + 500000) / 1000000 + (in15 * W15 + 500000) / 1000000;
    sum_0_8 <= (in16 * W16 + 500000) / 1000000 + (in17 * W17 + 500000) / 1000000;
    sum_0_9 <= (in18 * W18 + 500000) / 1000000 + (in19 * W19 + 500000) / 1000000;
    sum_0_10 <= (in20 * W20 + 500000) / 1000000 + (in21 * W21 + 500000) / 1000000;
    sum_0_11 <= (in22 * W22 + 500000) / 1000000 + (in23 * W23 + 500000) / 1000000;
    sum_0_12 <= (in24 * W24 + 500000) / 1000000 + (in25 * W25 + 500000) / 1000000;
    sum_0_13 <= (in26 * W26 + 500000) / 1000000 + (in27 * W27 + 500000) / 1000000;
    sum_0_14 <= (in28 * W28 + 500000) / 1000000 + (in29 * W29 + 500000) / 1000000;
    sum_0_15 <= (in30 * W30 + 500000) / 1000000 + (in31 * W31 + 500000) / 1000000;
    sum_0_16 <= (in32 * W32 + 500000) / 1000000 + (in33 * W33 + 500000) / 1000000;
    sum_0_17 <= (in34 * W34 + 500000) / 1000000 + (in35 * W35 + 500000) / 1000000;
    sum_0_18 <= (in36 * W36 + 500000) / 1000000 + (in37 * W37 + 500000) / 1000000;
    sum_0_19 <= (in38 * W38 + 500000) / 1000000 + (in39 * W39 + 500000) / 1000000;
    sum_0_20 <= (in40 * W40 + 500000) / 1000000 + (in41 * W41 + 500000) / 1000000;
    sum_0_21 <= (in42 * W42 + 500000) / 1000000 + (in43 * W43 + 500000) / 1000000;
    sum_0_22 <= (in44 * W44 + 500000) / 1000000 + (in45 * W45 + 500000) / 1000000;
    sum_0_23 <= (in46 * W46 + 500000) / 1000000 + (in47 * W47 + 500000) / 1000000;
    sum_0_24 <= (in48 * W48 + 500000) / 1000000 + (in49 * W49 + 500000) / 1000000;
    sum_0_25 <= (in50 * W50 + 500000) / 1000000 + (in51 * W51 + 500000) / 1000000;
    sum_0_26 <= (in52 * W52 + 500000) / 1000000 + (in53 * W53 + 500000) / 1000000;
    sum_0_27 <= (in54 * W54 + 500000) / 1000000 + (in55 * W55 + 500000) / 1000000;
    sum_0_28 <= (in56 * W56 + 500000) / 1000000 + (in57 * W57 + 500000) / 1000000;
    sum_0_29 <= (in58 * W58 + 500000) / 1000000 + (in59 * W59 + 500000) / 1000000;
    sum_0_30 <= (in60 * W60 + 500000) / 1000000 + (in61 * W61 + 500000) / 1000000;
    sum_0_31 <= (in62 * W62 + 500000) / 1000000 + (in63 * W63 + 500000) / 1000000 + BIAS;
    sum_1_0 <= sum_0_0 + sum_0_1;
    sum_1_1 <= sum_0_2 + sum_0_3;
    sum_1_2 <= sum_0_4 + sum_0_5;
    sum_1_3 <= sum_0_6 + sum_0_7;
    sum_1_4 <= sum_0_8 + sum_0_9;
    sum_1_5 <= sum_0_10 + sum_0_11;
    sum_1_6 <= sum_0_12 + sum_0_13;
    sum_1_7 <= sum_0_14 + sum_0_15;
    sum_1_8 <= sum_0_16 + sum_0_17;
    sum_1_9 <= sum_0_18 + sum_0_19;
    sum_1_10 <= sum_0_20 + sum_0_21;
    sum_1_11 <= sum_0_22 + sum_0_23;
    sum_1_12 <= sum_0_24 + sum_0_25;
    sum_1_13 <= sum_0_26 + sum_0_27;
    sum_1_14 <= sum_0_28 + sum_0_29;
    sum_1_15 <= sum_0_30 + sum_0_31;
    sum_2_0 <= sum_1_0 + sum_1_1;
    sum_2_1 <= sum_1_2 + sum_1_3;
    sum_2_2 <= sum_1_4 + sum_1_5;
    sum_2_3 <= sum_1_6 + sum_1_7;
    sum_2_4 <= sum_1_8 + sum_1_9;
    sum_2_5 <= sum_1_10 + sum_1_11;
    sum_2_6 <= sum_1_12 + sum_1_13;
    sum_2_7 <= sum_1_14 + sum_1_15;
    sum_3_0 <= sum_2_0 + sum_2_1;
    sum_3_1 <= sum_2_2 + sum_2_3;
    sum_3_2 <= sum_2_4 + sum_2_5;
    sum_3_3 <= sum_2_6 + sum_2_7;
    sum_4_0 <= sum_3_0 + sum_3_1;
    sum_4_1 <= sum_3_2 + sum_3_3;
    sum_5_0 <= sum_4_0 + sum_4_1;
    x <= sum_5_0;
    abs_x = x < 0 ? -x : x;
    if (abs_x >= 5000000) y = 1000000;
    else if (abs_x >= 2375000) y = 31250 * abs_x / 1000000 + 843750;
    else if (abs_x >= 1000000) y = 125000 * abs_x / 1000000 + 625000;
    else y = 250000 * abs_x / 1000000 + 500000;
    out = x < 0 ? 1000000 - y : y;
end

endmodule

module layer65in64out(clk, rst, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, out0, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13, out14, out15, out16, out17, out18, out19, out20, out21, out22, out23, out24, out25, out26, out27, out28, out29, out30, out31, out32, out33, out34, out35, out36, out37, out38, out39, out40, out41, out42, out43, out44, out45, out46, out47, out48, out49, out50, out51, out52, out53, out54, out55, out56, out57, out58, out59, out60, out61, out62, out63);

parameter signed BIAS0 = 0;
parameter signed BIAS1 = 0;
parameter signed BIAS2 = 0;
parameter signed BIAS3 = 0;
parameter signed BIAS4 = 0;
parameter signed BIAS5 = 0;
parameter signed BIAS6 = 0;
parameter signed BIAS7 = 0;
parameter signed BIAS8 = 0;
parameter signed BIAS9 = 0;
parameter signed BIAS10 = 0;
parameter signed BIAS11 = 0;
parameter signed BIAS12 = 0;
parameter signed BIAS13 = 0;
parameter signed BIAS14 = 0;
parameter signed BIAS15 = 0;
parameter signed BIAS16 = 0;
parameter signed BIAS17 = 0;
parameter signed BIAS18 = 0;
parameter signed BIAS19 = 0;
parameter signed BIAS20 = 0;
parameter signed BIAS21 = 0;
parameter signed BIAS22 = 0;
parameter signed BIAS23 = 0;
parameter signed BIAS24 = 0;
parameter signed BIAS25 = 0;
parameter signed BIAS26 = 0;
parameter signed BIAS27 = 0;
parameter signed BIAS28 = 0;
parameter signed BIAS29 = 0;
parameter signed BIAS30 = 0;
parameter signed BIAS31 = 0;
parameter signed BIAS32 = 0;
parameter signed BIAS33 = 0;
parameter signed BIAS34 = 0;
parameter signed BIAS35 = 0;
parameter signed BIAS36 = 0;
parameter signed BIAS37 = 0;
parameter signed BIAS38 = 0;
parameter signed BIAS39 = 0;
parameter signed BIAS40 = 0;
parameter signed BIAS41 = 0;
parameter signed BIAS42 = 0;
parameter signed BIAS43 = 0;
parameter signed BIAS44 = 0;
parameter signed BIAS45 = 0;
parameter signed BIAS46 = 0;
parameter signed BIAS47 = 0;
parameter signed BIAS48 = 0;
parameter signed BIAS49 = 0;
parameter signed BIAS50 = 0;
parameter signed BIAS51 = 0;
parameter signed BIAS52 = 0;
parameter signed BIAS53 = 0;
parameter signed BIAS54 = 0;
parameter signed BIAS55 = 0;
parameter signed BIAS56 = 0;
parameter signed BIAS57 = 0;
parameter signed BIAS58 = 0;
parameter signed BIAS59 = 0;
parameter signed BIAS60 = 0;
parameter signed BIAS61 = 0;
parameter signed BIAS62 = 0;
parameter signed BIAS63 = 0;
parameter signed W0TO0 = 0;
parameter signed W0TO1 = 0;
parameter signed W0TO2 = 0;
parameter signed W0TO3 = 0;
parameter signed W0TO4 = 0;
parameter signed W0TO5 = 0;
parameter signed W0TO6 = 0;
parameter signed W0TO7 = 0;
parameter signed W0TO8 = 0;
parameter signed W0TO9 = 0;
parameter signed W0TO10 = 0;
parameter signed W0TO11 = 0;
parameter signed W0TO12 = 0;
parameter signed W0TO13 = 0;
parameter signed W0TO14 = 0;
parameter signed W0TO15 = 0;
parameter signed W0TO16 = 0;
parameter signed W0TO17 = 0;
parameter signed W0TO18 = 0;
parameter signed W0TO19 = 0;
parameter signed W0TO20 = 0;
parameter signed W0TO21 = 0;
parameter signed W0TO22 = 0;
parameter signed W0TO23 = 0;
parameter signed W0TO24 = 0;
parameter signed W0TO25 = 0;
parameter signed W0TO26 = 0;
parameter signed W0TO27 = 0;
parameter signed W0TO28 = 0;
parameter signed W0TO29 = 0;
parameter signed W0TO30 = 0;
parameter signed W0TO31 = 0;
parameter signed W0TO32 = 0;
parameter signed W0TO33 = 0;
parameter signed W0TO34 = 0;
parameter signed W0TO35 = 0;
parameter signed W0TO36 = 0;
parameter signed W0TO37 = 0;
parameter signed W0TO38 = 0;
parameter signed W0TO39 = 0;
parameter signed W0TO40 = 0;
parameter signed W0TO41 = 0;
parameter signed W0TO42 = 0;
parameter signed W0TO43 = 0;
parameter signed W0TO44 = 0;
parameter signed W0TO45 = 0;
parameter signed W0TO46 = 0;
parameter signed W0TO47 = 0;
parameter signed W0TO48 = 0;
parameter signed W0TO49 = 0;
parameter signed W0TO50 = 0;
parameter signed W0TO51 = 0;
parameter signed W0TO52 = 0;
parameter signed W0TO53 = 0;
parameter signed W0TO54 = 0;
parameter signed W0TO55 = 0;
parameter signed W0TO56 = 0;
parameter signed W0TO57 = 0;
parameter signed W0TO58 = 0;
parameter signed W0TO59 = 0;
parameter signed W0TO60 = 0;
parameter signed W0TO61 = 0;
parameter signed W0TO62 = 0;
parameter signed W0TO63 = 0;
parameter signed W1TO0 = 0;
parameter signed W1TO1 = 0;
parameter signed W1TO2 = 0;
parameter signed W1TO3 = 0;
parameter signed W1TO4 = 0;
parameter signed W1TO5 = 0;
parameter signed W1TO6 = 0;
parameter signed W1TO7 = 0;
parameter signed W1TO8 = 0;
parameter signed W1TO9 = 0;
parameter signed W1TO10 = 0;
parameter signed W1TO11 = 0;
parameter signed W1TO12 = 0;
parameter signed W1TO13 = 0;
parameter signed W1TO14 = 0;
parameter signed W1TO15 = 0;
parameter signed W1TO16 = 0;
parameter signed W1TO17 = 0;
parameter signed W1TO18 = 0;
parameter signed W1TO19 = 0;
parameter signed W1TO20 = 0;
parameter signed W1TO21 = 0;
parameter signed W1TO22 = 0;
parameter signed W1TO23 = 0;
parameter signed W1TO24 = 0;
parameter signed W1TO25 = 0;
parameter signed W1TO26 = 0;
parameter signed W1TO27 = 0;
parameter signed W1TO28 = 0;
parameter signed W1TO29 = 0;
parameter signed W1TO30 = 0;
parameter signed W1TO31 = 0;
parameter signed W1TO32 = 0;
parameter signed W1TO33 = 0;
parameter signed W1TO34 = 0;
parameter signed W1TO35 = 0;
parameter signed W1TO36 = 0;
parameter signed W1TO37 = 0;
parameter signed W1TO38 = 0;
parameter signed W1TO39 = 0;
parameter signed W1TO40 = 0;
parameter signed W1TO41 = 0;
parameter signed W1TO42 = 0;
parameter signed W1TO43 = 0;
parameter signed W1TO44 = 0;
parameter signed W1TO45 = 0;
parameter signed W1TO46 = 0;
parameter signed W1TO47 = 0;
parameter signed W1TO48 = 0;
parameter signed W1TO49 = 0;
parameter signed W1TO50 = 0;
parameter signed W1TO51 = 0;
parameter signed W1TO52 = 0;
parameter signed W1TO53 = 0;
parameter signed W1TO54 = 0;
parameter signed W1TO55 = 0;
parameter signed W1TO56 = 0;
parameter signed W1TO57 = 0;
parameter signed W1TO58 = 0;
parameter signed W1TO59 = 0;
parameter signed W1TO60 = 0;
parameter signed W1TO61 = 0;
parameter signed W1TO62 = 0;
parameter signed W1TO63 = 0;
parameter signed W2TO0 = 0;
parameter signed W2TO1 = 0;
parameter signed W2TO2 = 0;
parameter signed W2TO3 = 0;
parameter signed W2TO4 = 0;
parameter signed W2TO5 = 0;
parameter signed W2TO6 = 0;
parameter signed W2TO7 = 0;
parameter signed W2TO8 = 0;
parameter signed W2TO9 = 0;
parameter signed W2TO10 = 0;
parameter signed W2TO11 = 0;
parameter signed W2TO12 = 0;
parameter signed W2TO13 = 0;
parameter signed W2TO14 = 0;
parameter signed W2TO15 = 0;
parameter signed W2TO16 = 0;
parameter signed W2TO17 = 0;
parameter signed W2TO18 = 0;
parameter signed W2TO19 = 0;
parameter signed W2TO20 = 0;
parameter signed W2TO21 = 0;
parameter signed W2TO22 = 0;
parameter signed W2TO23 = 0;
parameter signed W2TO24 = 0;
parameter signed W2TO25 = 0;
parameter signed W2TO26 = 0;
parameter signed W2TO27 = 0;
parameter signed W2TO28 = 0;
parameter signed W2TO29 = 0;
parameter signed W2TO30 = 0;
parameter signed W2TO31 = 0;
parameter signed W2TO32 = 0;
parameter signed W2TO33 = 0;
parameter signed W2TO34 = 0;
parameter signed W2TO35 = 0;
parameter signed W2TO36 = 0;
parameter signed W2TO37 = 0;
parameter signed W2TO38 = 0;
parameter signed W2TO39 = 0;
parameter signed W2TO40 = 0;
parameter signed W2TO41 = 0;
parameter signed W2TO42 = 0;
parameter signed W2TO43 = 0;
parameter signed W2TO44 = 0;
parameter signed W2TO45 = 0;
parameter signed W2TO46 = 0;
parameter signed W2TO47 = 0;
parameter signed W2TO48 = 0;
parameter signed W2TO49 = 0;
parameter signed W2TO50 = 0;
parameter signed W2TO51 = 0;
parameter signed W2TO52 = 0;
parameter signed W2TO53 = 0;
parameter signed W2TO54 = 0;
parameter signed W2TO55 = 0;
parameter signed W2TO56 = 0;
parameter signed W2TO57 = 0;
parameter signed W2TO58 = 0;
parameter signed W2TO59 = 0;
parameter signed W2TO60 = 0;
parameter signed W2TO61 = 0;
parameter signed W2TO62 = 0;
parameter signed W2TO63 = 0;
parameter signed W3TO0 = 0;
parameter signed W3TO1 = 0;
parameter signed W3TO2 = 0;
parameter signed W3TO3 = 0;
parameter signed W3TO4 = 0;
parameter signed W3TO5 = 0;
parameter signed W3TO6 = 0;
parameter signed W3TO7 = 0;
parameter signed W3TO8 = 0;
parameter signed W3TO9 = 0;
parameter signed W3TO10 = 0;
parameter signed W3TO11 = 0;
parameter signed W3TO12 = 0;
parameter signed W3TO13 = 0;
parameter signed W3TO14 = 0;
parameter signed W3TO15 = 0;
parameter signed W3TO16 = 0;
parameter signed W3TO17 = 0;
parameter signed W3TO18 = 0;
parameter signed W3TO19 = 0;
parameter signed W3TO20 = 0;
parameter signed W3TO21 = 0;
parameter signed W3TO22 = 0;
parameter signed W3TO23 = 0;
parameter signed W3TO24 = 0;
parameter signed W3TO25 = 0;
parameter signed W3TO26 = 0;
parameter signed W3TO27 = 0;
parameter signed W3TO28 = 0;
parameter signed W3TO29 = 0;
parameter signed W3TO30 = 0;
parameter signed W3TO31 = 0;
parameter signed W3TO32 = 0;
parameter signed W3TO33 = 0;
parameter signed W3TO34 = 0;
parameter signed W3TO35 = 0;
parameter signed W3TO36 = 0;
parameter signed W3TO37 = 0;
parameter signed W3TO38 = 0;
parameter signed W3TO39 = 0;
parameter signed W3TO40 = 0;
parameter signed W3TO41 = 0;
parameter signed W3TO42 = 0;
parameter signed W3TO43 = 0;
parameter signed W3TO44 = 0;
parameter signed W3TO45 = 0;
parameter signed W3TO46 = 0;
parameter signed W3TO47 = 0;
parameter signed W3TO48 = 0;
parameter signed W3TO49 = 0;
parameter signed W3TO50 = 0;
parameter signed W3TO51 = 0;
parameter signed W3TO52 = 0;
parameter signed W3TO53 = 0;
parameter signed W3TO54 = 0;
parameter signed W3TO55 = 0;
parameter signed W3TO56 = 0;
parameter signed W3TO57 = 0;
parameter signed W3TO58 = 0;
parameter signed W3TO59 = 0;
parameter signed W3TO60 = 0;
parameter signed W3TO61 = 0;
parameter signed W3TO62 = 0;
parameter signed W3TO63 = 0;
parameter signed W4TO0 = 0;
parameter signed W4TO1 = 0;
parameter signed W4TO2 = 0;
parameter signed W4TO3 = 0;
parameter signed W4TO4 = 0;
parameter signed W4TO5 = 0;
parameter signed W4TO6 = 0;
parameter signed W4TO7 = 0;
parameter signed W4TO8 = 0;
parameter signed W4TO9 = 0;
parameter signed W4TO10 = 0;
parameter signed W4TO11 = 0;
parameter signed W4TO12 = 0;
parameter signed W4TO13 = 0;
parameter signed W4TO14 = 0;
parameter signed W4TO15 = 0;
parameter signed W4TO16 = 0;
parameter signed W4TO17 = 0;
parameter signed W4TO18 = 0;
parameter signed W4TO19 = 0;
parameter signed W4TO20 = 0;
parameter signed W4TO21 = 0;
parameter signed W4TO22 = 0;
parameter signed W4TO23 = 0;
parameter signed W4TO24 = 0;
parameter signed W4TO25 = 0;
parameter signed W4TO26 = 0;
parameter signed W4TO27 = 0;
parameter signed W4TO28 = 0;
parameter signed W4TO29 = 0;
parameter signed W4TO30 = 0;
parameter signed W4TO31 = 0;
parameter signed W4TO32 = 0;
parameter signed W4TO33 = 0;
parameter signed W4TO34 = 0;
parameter signed W4TO35 = 0;
parameter signed W4TO36 = 0;
parameter signed W4TO37 = 0;
parameter signed W4TO38 = 0;
parameter signed W4TO39 = 0;
parameter signed W4TO40 = 0;
parameter signed W4TO41 = 0;
parameter signed W4TO42 = 0;
parameter signed W4TO43 = 0;
parameter signed W4TO44 = 0;
parameter signed W4TO45 = 0;
parameter signed W4TO46 = 0;
parameter signed W4TO47 = 0;
parameter signed W4TO48 = 0;
parameter signed W4TO49 = 0;
parameter signed W4TO50 = 0;
parameter signed W4TO51 = 0;
parameter signed W4TO52 = 0;
parameter signed W4TO53 = 0;
parameter signed W4TO54 = 0;
parameter signed W4TO55 = 0;
parameter signed W4TO56 = 0;
parameter signed W4TO57 = 0;
parameter signed W4TO58 = 0;
parameter signed W4TO59 = 0;
parameter signed W4TO60 = 0;
parameter signed W4TO61 = 0;
parameter signed W4TO62 = 0;
parameter signed W4TO63 = 0;
parameter signed W5TO0 = 0;
parameter signed W5TO1 = 0;
parameter signed W5TO2 = 0;
parameter signed W5TO3 = 0;
parameter signed W5TO4 = 0;
parameter signed W5TO5 = 0;
parameter signed W5TO6 = 0;
parameter signed W5TO7 = 0;
parameter signed W5TO8 = 0;
parameter signed W5TO9 = 0;
parameter signed W5TO10 = 0;
parameter signed W5TO11 = 0;
parameter signed W5TO12 = 0;
parameter signed W5TO13 = 0;
parameter signed W5TO14 = 0;
parameter signed W5TO15 = 0;
parameter signed W5TO16 = 0;
parameter signed W5TO17 = 0;
parameter signed W5TO18 = 0;
parameter signed W5TO19 = 0;
parameter signed W5TO20 = 0;
parameter signed W5TO21 = 0;
parameter signed W5TO22 = 0;
parameter signed W5TO23 = 0;
parameter signed W5TO24 = 0;
parameter signed W5TO25 = 0;
parameter signed W5TO26 = 0;
parameter signed W5TO27 = 0;
parameter signed W5TO28 = 0;
parameter signed W5TO29 = 0;
parameter signed W5TO30 = 0;
parameter signed W5TO31 = 0;
parameter signed W5TO32 = 0;
parameter signed W5TO33 = 0;
parameter signed W5TO34 = 0;
parameter signed W5TO35 = 0;
parameter signed W5TO36 = 0;
parameter signed W5TO37 = 0;
parameter signed W5TO38 = 0;
parameter signed W5TO39 = 0;
parameter signed W5TO40 = 0;
parameter signed W5TO41 = 0;
parameter signed W5TO42 = 0;
parameter signed W5TO43 = 0;
parameter signed W5TO44 = 0;
parameter signed W5TO45 = 0;
parameter signed W5TO46 = 0;
parameter signed W5TO47 = 0;
parameter signed W5TO48 = 0;
parameter signed W5TO49 = 0;
parameter signed W5TO50 = 0;
parameter signed W5TO51 = 0;
parameter signed W5TO52 = 0;
parameter signed W5TO53 = 0;
parameter signed W5TO54 = 0;
parameter signed W5TO55 = 0;
parameter signed W5TO56 = 0;
parameter signed W5TO57 = 0;
parameter signed W5TO58 = 0;
parameter signed W5TO59 = 0;
parameter signed W5TO60 = 0;
parameter signed W5TO61 = 0;
parameter signed W5TO62 = 0;
parameter signed W5TO63 = 0;
parameter signed W6TO0 = 0;
parameter signed W6TO1 = 0;
parameter signed W6TO2 = 0;
parameter signed W6TO3 = 0;
parameter signed W6TO4 = 0;
parameter signed W6TO5 = 0;
parameter signed W6TO6 = 0;
parameter signed W6TO7 = 0;
parameter signed W6TO8 = 0;
parameter signed W6TO9 = 0;
parameter signed W6TO10 = 0;
parameter signed W6TO11 = 0;
parameter signed W6TO12 = 0;
parameter signed W6TO13 = 0;
parameter signed W6TO14 = 0;
parameter signed W6TO15 = 0;
parameter signed W6TO16 = 0;
parameter signed W6TO17 = 0;
parameter signed W6TO18 = 0;
parameter signed W6TO19 = 0;
parameter signed W6TO20 = 0;
parameter signed W6TO21 = 0;
parameter signed W6TO22 = 0;
parameter signed W6TO23 = 0;
parameter signed W6TO24 = 0;
parameter signed W6TO25 = 0;
parameter signed W6TO26 = 0;
parameter signed W6TO27 = 0;
parameter signed W6TO28 = 0;
parameter signed W6TO29 = 0;
parameter signed W6TO30 = 0;
parameter signed W6TO31 = 0;
parameter signed W6TO32 = 0;
parameter signed W6TO33 = 0;
parameter signed W6TO34 = 0;
parameter signed W6TO35 = 0;
parameter signed W6TO36 = 0;
parameter signed W6TO37 = 0;
parameter signed W6TO38 = 0;
parameter signed W6TO39 = 0;
parameter signed W6TO40 = 0;
parameter signed W6TO41 = 0;
parameter signed W6TO42 = 0;
parameter signed W6TO43 = 0;
parameter signed W6TO44 = 0;
parameter signed W6TO45 = 0;
parameter signed W6TO46 = 0;
parameter signed W6TO47 = 0;
parameter signed W6TO48 = 0;
parameter signed W6TO49 = 0;
parameter signed W6TO50 = 0;
parameter signed W6TO51 = 0;
parameter signed W6TO52 = 0;
parameter signed W6TO53 = 0;
parameter signed W6TO54 = 0;
parameter signed W6TO55 = 0;
parameter signed W6TO56 = 0;
parameter signed W6TO57 = 0;
parameter signed W6TO58 = 0;
parameter signed W6TO59 = 0;
parameter signed W6TO60 = 0;
parameter signed W6TO61 = 0;
parameter signed W6TO62 = 0;
parameter signed W6TO63 = 0;
parameter signed W7TO0 = 0;
parameter signed W7TO1 = 0;
parameter signed W7TO2 = 0;
parameter signed W7TO3 = 0;
parameter signed W7TO4 = 0;
parameter signed W7TO5 = 0;
parameter signed W7TO6 = 0;
parameter signed W7TO7 = 0;
parameter signed W7TO8 = 0;
parameter signed W7TO9 = 0;
parameter signed W7TO10 = 0;
parameter signed W7TO11 = 0;
parameter signed W7TO12 = 0;
parameter signed W7TO13 = 0;
parameter signed W7TO14 = 0;
parameter signed W7TO15 = 0;
parameter signed W7TO16 = 0;
parameter signed W7TO17 = 0;
parameter signed W7TO18 = 0;
parameter signed W7TO19 = 0;
parameter signed W7TO20 = 0;
parameter signed W7TO21 = 0;
parameter signed W7TO22 = 0;
parameter signed W7TO23 = 0;
parameter signed W7TO24 = 0;
parameter signed W7TO25 = 0;
parameter signed W7TO26 = 0;
parameter signed W7TO27 = 0;
parameter signed W7TO28 = 0;
parameter signed W7TO29 = 0;
parameter signed W7TO30 = 0;
parameter signed W7TO31 = 0;
parameter signed W7TO32 = 0;
parameter signed W7TO33 = 0;
parameter signed W7TO34 = 0;
parameter signed W7TO35 = 0;
parameter signed W7TO36 = 0;
parameter signed W7TO37 = 0;
parameter signed W7TO38 = 0;
parameter signed W7TO39 = 0;
parameter signed W7TO40 = 0;
parameter signed W7TO41 = 0;
parameter signed W7TO42 = 0;
parameter signed W7TO43 = 0;
parameter signed W7TO44 = 0;
parameter signed W7TO45 = 0;
parameter signed W7TO46 = 0;
parameter signed W7TO47 = 0;
parameter signed W7TO48 = 0;
parameter signed W7TO49 = 0;
parameter signed W7TO50 = 0;
parameter signed W7TO51 = 0;
parameter signed W7TO52 = 0;
parameter signed W7TO53 = 0;
parameter signed W7TO54 = 0;
parameter signed W7TO55 = 0;
parameter signed W7TO56 = 0;
parameter signed W7TO57 = 0;
parameter signed W7TO58 = 0;
parameter signed W7TO59 = 0;
parameter signed W7TO60 = 0;
parameter signed W7TO61 = 0;
parameter signed W7TO62 = 0;
parameter signed W7TO63 = 0;
parameter signed W8TO0 = 0;
parameter signed W8TO1 = 0;
parameter signed W8TO2 = 0;
parameter signed W8TO3 = 0;
parameter signed W8TO4 = 0;
parameter signed W8TO5 = 0;
parameter signed W8TO6 = 0;
parameter signed W8TO7 = 0;
parameter signed W8TO8 = 0;
parameter signed W8TO9 = 0;
parameter signed W8TO10 = 0;
parameter signed W8TO11 = 0;
parameter signed W8TO12 = 0;
parameter signed W8TO13 = 0;
parameter signed W8TO14 = 0;
parameter signed W8TO15 = 0;
parameter signed W8TO16 = 0;
parameter signed W8TO17 = 0;
parameter signed W8TO18 = 0;
parameter signed W8TO19 = 0;
parameter signed W8TO20 = 0;
parameter signed W8TO21 = 0;
parameter signed W8TO22 = 0;
parameter signed W8TO23 = 0;
parameter signed W8TO24 = 0;
parameter signed W8TO25 = 0;
parameter signed W8TO26 = 0;
parameter signed W8TO27 = 0;
parameter signed W8TO28 = 0;
parameter signed W8TO29 = 0;
parameter signed W8TO30 = 0;
parameter signed W8TO31 = 0;
parameter signed W8TO32 = 0;
parameter signed W8TO33 = 0;
parameter signed W8TO34 = 0;
parameter signed W8TO35 = 0;
parameter signed W8TO36 = 0;
parameter signed W8TO37 = 0;
parameter signed W8TO38 = 0;
parameter signed W8TO39 = 0;
parameter signed W8TO40 = 0;
parameter signed W8TO41 = 0;
parameter signed W8TO42 = 0;
parameter signed W8TO43 = 0;
parameter signed W8TO44 = 0;
parameter signed W8TO45 = 0;
parameter signed W8TO46 = 0;
parameter signed W8TO47 = 0;
parameter signed W8TO48 = 0;
parameter signed W8TO49 = 0;
parameter signed W8TO50 = 0;
parameter signed W8TO51 = 0;
parameter signed W8TO52 = 0;
parameter signed W8TO53 = 0;
parameter signed W8TO54 = 0;
parameter signed W8TO55 = 0;
parameter signed W8TO56 = 0;
parameter signed W8TO57 = 0;
parameter signed W8TO58 = 0;
parameter signed W8TO59 = 0;
parameter signed W8TO60 = 0;
parameter signed W8TO61 = 0;
parameter signed W8TO62 = 0;
parameter signed W8TO63 = 0;
parameter signed W9TO0 = 0;
parameter signed W9TO1 = 0;
parameter signed W9TO2 = 0;
parameter signed W9TO3 = 0;
parameter signed W9TO4 = 0;
parameter signed W9TO5 = 0;
parameter signed W9TO6 = 0;
parameter signed W9TO7 = 0;
parameter signed W9TO8 = 0;
parameter signed W9TO9 = 0;
parameter signed W9TO10 = 0;
parameter signed W9TO11 = 0;
parameter signed W9TO12 = 0;
parameter signed W9TO13 = 0;
parameter signed W9TO14 = 0;
parameter signed W9TO15 = 0;
parameter signed W9TO16 = 0;
parameter signed W9TO17 = 0;
parameter signed W9TO18 = 0;
parameter signed W9TO19 = 0;
parameter signed W9TO20 = 0;
parameter signed W9TO21 = 0;
parameter signed W9TO22 = 0;
parameter signed W9TO23 = 0;
parameter signed W9TO24 = 0;
parameter signed W9TO25 = 0;
parameter signed W9TO26 = 0;
parameter signed W9TO27 = 0;
parameter signed W9TO28 = 0;
parameter signed W9TO29 = 0;
parameter signed W9TO30 = 0;
parameter signed W9TO31 = 0;
parameter signed W9TO32 = 0;
parameter signed W9TO33 = 0;
parameter signed W9TO34 = 0;
parameter signed W9TO35 = 0;
parameter signed W9TO36 = 0;
parameter signed W9TO37 = 0;
parameter signed W9TO38 = 0;
parameter signed W9TO39 = 0;
parameter signed W9TO40 = 0;
parameter signed W9TO41 = 0;
parameter signed W9TO42 = 0;
parameter signed W9TO43 = 0;
parameter signed W9TO44 = 0;
parameter signed W9TO45 = 0;
parameter signed W9TO46 = 0;
parameter signed W9TO47 = 0;
parameter signed W9TO48 = 0;
parameter signed W9TO49 = 0;
parameter signed W9TO50 = 0;
parameter signed W9TO51 = 0;
parameter signed W9TO52 = 0;
parameter signed W9TO53 = 0;
parameter signed W9TO54 = 0;
parameter signed W9TO55 = 0;
parameter signed W9TO56 = 0;
parameter signed W9TO57 = 0;
parameter signed W9TO58 = 0;
parameter signed W9TO59 = 0;
parameter signed W9TO60 = 0;
parameter signed W9TO61 = 0;
parameter signed W9TO62 = 0;
parameter signed W9TO63 = 0;
parameter signed W10TO0 = 0;
parameter signed W10TO1 = 0;
parameter signed W10TO2 = 0;
parameter signed W10TO3 = 0;
parameter signed W10TO4 = 0;
parameter signed W10TO5 = 0;
parameter signed W10TO6 = 0;
parameter signed W10TO7 = 0;
parameter signed W10TO8 = 0;
parameter signed W10TO9 = 0;
parameter signed W10TO10 = 0;
parameter signed W10TO11 = 0;
parameter signed W10TO12 = 0;
parameter signed W10TO13 = 0;
parameter signed W10TO14 = 0;
parameter signed W10TO15 = 0;
parameter signed W10TO16 = 0;
parameter signed W10TO17 = 0;
parameter signed W10TO18 = 0;
parameter signed W10TO19 = 0;
parameter signed W10TO20 = 0;
parameter signed W10TO21 = 0;
parameter signed W10TO22 = 0;
parameter signed W10TO23 = 0;
parameter signed W10TO24 = 0;
parameter signed W10TO25 = 0;
parameter signed W10TO26 = 0;
parameter signed W10TO27 = 0;
parameter signed W10TO28 = 0;
parameter signed W10TO29 = 0;
parameter signed W10TO30 = 0;
parameter signed W10TO31 = 0;
parameter signed W10TO32 = 0;
parameter signed W10TO33 = 0;
parameter signed W10TO34 = 0;
parameter signed W10TO35 = 0;
parameter signed W10TO36 = 0;
parameter signed W10TO37 = 0;
parameter signed W10TO38 = 0;
parameter signed W10TO39 = 0;
parameter signed W10TO40 = 0;
parameter signed W10TO41 = 0;
parameter signed W10TO42 = 0;
parameter signed W10TO43 = 0;
parameter signed W10TO44 = 0;
parameter signed W10TO45 = 0;
parameter signed W10TO46 = 0;
parameter signed W10TO47 = 0;
parameter signed W10TO48 = 0;
parameter signed W10TO49 = 0;
parameter signed W10TO50 = 0;
parameter signed W10TO51 = 0;
parameter signed W10TO52 = 0;
parameter signed W10TO53 = 0;
parameter signed W10TO54 = 0;
parameter signed W10TO55 = 0;
parameter signed W10TO56 = 0;
parameter signed W10TO57 = 0;
parameter signed W10TO58 = 0;
parameter signed W10TO59 = 0;
parameter signed W10TO60 = 0;
parameter signed W10TO61 = 0;
parameter signed W10TO62 = 0;
parameter signed W10TO63 = 0;
parameter signed W11TO0 = 0;
parameter signed W11TO1 = 0;
parameter signed W11TO2 = 0;
parameter signed W11TO3 = 0;
parameter signed W11TO4 = 0;
parameter signed W11TO5 = 0;
parameter signed W11TO6 = 0;
parameter signed W11TO7 = 0;
parameter signed W11TO8 = 0;
parameter signed W11TO9 = 0;
parameter signed W11TO10 = 0;
parameter signed W11TO11 = 0;
parameter signed W11TO12 = 0;
parameter signed W11TO13 = 0;
parameter signed W11TO14 = 0;
parameter signed W11TO15 = 0;
parameter signed W11TO16 = 0;
parameter signed W11TO17 = 0;
parameter signed W11TO18 = 0;
parameter signed W11TO19 = 0;
parameter signed W11TO20 = 0;
parameter signed W11TO21 = 0;
parameter signed W11TO22 = 0;
parameter signed W11TO23 = 0;
parameter signed W11TO24 = 0;
parameter signed W11TO25 = 0;
parameter signed W11TO26 = 0;
parameter signed W11TO27 = 0;
parameter signed W11TO28 = 0;
parameter signed W11TO29 = 0;
parameter signed W11TO30 = 0;
parameter signed W11TO31 = 0;
parameter signed W11TO32 = 0;
parameter signed W11TO33 = 0;
parameter signed W11TO34 = 0;
parameter signed W11TO35 = 0;
parameter signed W11TO36 = 0;
parameter signed W11TO37 = 0;
parameter signed W11TO38 = 0;
parameter signed W11TO39 = 0;
parameter signed W11TO40 = 0;
parameter signed W11TO41 = 0;
parameter signed W11TO42 = 0;
parameter signed W11TO43 = 0;
parameter signed W11TO44 = 0;
parameter signed W11TO45 = 0;
parameter signed W11TO46 = 0;
parameter signed W11TO47 = 0;
parameter signed W11TO48 = 0;
parameter signed W11TO49 = 0;
parameter signed W11TO50 = 0;
parameter signed W11TO51 = 0;
parameter signed W11TO52 = 0;
parameter signed W11TO53 = 0;
parameter signed W11TO54 = 0;
parameter signed W11TO55 = 0;
parameter signed W11TO56 = 0;
parameter signed W11TO57 = 0;
parameter signed W11TO58 = 0;
parameter signed W11TO59 = 0;
parameter signed W11TO60 = 0;
parameter signed W11TO61 = 0;
parameter signed W11TO62 = 0;
parameter signed W11TO63 = 0;
parameter signed W12TO0 = 0;
parameter signed W12TO1 = 0;
parameter signed W12TO2 = 0;
parameter signed W12TO3 = 0;
parameter signed W12TO4 = 0;
parameter signed W12TO5 = 0;
parameter signed W12TO6 = 0;
parameter signed W12TO7 = 0;
parameter signed W12TO8 = 0;
parameter signed W12TO9 = 0;
parameter signed W12TO10 = 0;
parameter signed W12TO11 = 0;
parameter signed W12TO12 = 0;
parameter signed W12TO13 = 0;
parameter signed W12TO14 = 0;
parameter signed W12TO15 = 0;
parameter signed W12TO16 = 0;
parameter signed W12TO17 = 0;
parameter signed W12TO18 = 0;
parameter signed W12TO19 = 0;
parameter signed W12TO20 = 0;
parameter signed W12TO21 = 0;
parameter signed W12TO22 = 0;
parameter signed W12TO23 = 0;
parameter signed W12TO24 = 0;
parameter signed W12TO25 = 0;
parameter signed W12TO26 = 0;
parameter signed W12TO27 = 0;
parameter signed W12TO28 = 0;
parameter signed W12TO29 = 0;
parameter signed W12TO30 = 0;
parameter signed W12TO31 = 0;
parameter signed W12TO32 = 0;
parameter signed W12TO33 = 0;
parameter signed W12TO34 = 0;
parameter signed W12TO35 = 0;
parameter signed W12TO36 = 0;
parameter signed W12TO37 = 0;
parameter signed W12TO38 = 0;
parameter signed W12TO39 = 0;
parameter signed W12TO40 = 0;
parameter signed W12TO41 = 0;
parameter signed W12TO42 = 0;
parameter signed W12TO43 = 0;
parameter signed W12TO44 = 0;
parameter signed W12TO45 = 0;
parameter signed W12TO46 = 0;
parameter signed W12TO47 = 0;
parameter signed W12TO48 = 0;
parameter signed W12TO49 = 0;
parameter signed W12TO50 = 0;
parameter signed W12TO51 = 0;
parameter signed W12TO52 = 0;
parameter signed W12TO53 = 0;
parameter signed W12TO54 = 0;
parameter signed W12TO55 = 0;
parameter signed W12TO56 = 0;
parameter signed W12TO57 = 0;
parameter signed W12TO58 = 0;
parameter signed W12TO59 = 0;
parameter signed W12TO60 = 0;
parameter signed W12TO61 = 0;
parameter signed W12TO62 = 0;
parameter signed W12TO63 = 0;
parameter signed W13TO0 = 0;
parameter signed W13TO1 = 0;
parameter signed W13TO2 = 0;
parameter signed W13TO3 = 0;
parameter signed W13TO4 = 0;
parameter signed W13TO5 = 0;
parameter signed W13TO6 = 0;
parameter signed W13TO7 = 0;
parameter signed W13TO8 = 0;
parameter signed W13TO9 = 0;
parameter signed W13TO10 = 0;
parameter signed W13TO11 = 0;
parameter signed W13TO12 = 0;
parameter signed W13TO13 = 0;
parameter signed W13TO14 = 0;
parameter signed W13TO15 = 0;
parameter signed W13TO16 = 0;
parameter signed W13TO17 = 0;
parameter signed W13TO18 = 0;
parameter signed W13TO19 = 0;
parameter signed W13TO20 = 0;
parameter signed W13TO21 = 0;
parameter signed W13TO22 = 0;
parameter signed W13TO23 = 0;
parameter signed W13TO24 = 0;
parameter signed W13TO25 = 0;
parameter signed W13TO26 = 0;
parameter signed W13TO27 = 0;
parameter signed W13TO28 = 0;
parameter signed W13TO29 = 0;
parameter signed W13TO30 = 0;
parameter signed W13TO31 = 0;
parameter signed W13TO32 = 0;
parameter signed W13TO33 = 0;
parameter signed W13TO34 = 0;
parameter signed W13TO35 = 0;
parameter signed W13TO36 = 0;
parameter signed W13TO37 = 0;
parameter signed W13TO38 = 0;
parameter signed W13TO39 = 0;
parameter signed W13TO40 = 0;
parameter signed W13TO41 = 0;
parameter signed W13TO42 = 0;
parameter signed W13TO43 = 0;
parameter signed W13TO44 = 0;
parameter signed W13TO45 = 0;
parameter signed W13TO46 = 0;
parameter signed W13TO47 = 0;
parameter signed W13TO48 = 0;
parameter signed W13TO49 = 0;
parameter signed W13TO50 = 0;
parameter signed W13TO51 = 0;
parameter signed W13TO52 = 0;
parameter signed W13TO53 = 0;
parameter signed W13TO54 = 0;
parameter signed W13TO55 = 0;
parameter signed W13TO56 = 0;
parameter signed W13TO57 = 0;
parameter signed W13TO58 = 0;
parameter signed W13TO59 = 0;
parameter signed W13TO60 = 0;
parameter signed W13TO61 = 0;
parameter signed W13TO62 = 0;
parameter signed W13TO63 = 0;
parameter signed W14TO0 = 0;
parameter signed W14TO1 = 0;
parameter signed W14TO2 = 0;
parameter signed W14TO3 = 0;
parameter signed W14TO4 = 0;
parameter signed W14TO5 = 0;
parameter signed W14TO6 = 0;
parameter signed W14TO7 = 0;
parameter signed W14TO8 = 0;
parameter signed W14TO9 = 0;
parameter signed W14TO10 = 0;
parameter signed W14TO11 = 0;
parameter signed W14TO12 = 0;
parameter signed W14TO13 = 0;
parameter signed W14TO14 = 0;
parameter signed W14TO15 = 0;
parameter signed W14TO16 = 0;
parameter signed W14TO17 = 0;
parameter signed W14TO18 = 0;
parameter signed W14TO19 = 0;
parameter signed W14TO20 = 0;
parameter signed W14TO21 = 0;
parameter signed W14TO22 = 0;
parameter signed W14TO23 = 0;
parameter signed W14TO24 = 0;
parameter signed W14TO25 = 0;
parameter signed W14TO26 = 0;
parameter signed W14TO27 = 0;
parameter signed W14TO28 = 0;
parameter signed W14TO29 = 0;
parameter signed W14TO30 = 0;
parameter signed W14TO31 = 0;
parameter signed W14TO32 = 0;
parameter signed W14TO33 = 0;
parameter signed W14TO34 = 0;
parameter signed W14TO35 = 0;
parameter signed W14TO36 = 0;
parameter signed W14TO37 = 0;
parameter signed W14TO38 = 0;
parameter signed W14TO39 = 0;
parameter signed W14TO40 = 0;
parameter signed W14TO41 = 0;
parameter signed W14TO42 = 0;
parameter signed W14TO43 = 0;
parameter signed W14TO44 = 0;
parameter signed W14TO45 = 0;
parameter signed W14TO46 = 0;
parameter signed W14TO47 = 0;
parameter signed W14TO48 = 0;
parameter signed W14TO49 = 0;
parameter signed W14TO50 = 0;
parameter signed W14TO51 = 0;
parameter signed W14TO52 = 0;
parameter signed W14TO53 = 0;
parameter signed W14TO54 = 0;
parameter signed W14TO55 = 0;
parameter signed W14TO56 = 0;
parameter signed W14TO57 = 0;
parameter signed W14TO58 = 0;
parameter signed W14TO59 = 0;
parameter signed W14TO60 = 0;
parameter signed W14TO61 = 0;
parameter signed W14TO62 = 0;
parameter signed W14TO63 = 0;
parameter signed W15TO0 = 0;
parameter signed W15TO1 = 0;
parameter signed W15TO2 = 0;
parameter signed W15TO3 = 0;
parameter signed W15TO4 = 0;
parameter signed W15TO5 = 0;
parameter signed W15TO6 = 0;
parameter signed W15TO7 = 0;
parameter signed W15TO8 = 0;
parameter signed W15TO9 = 0;
parameter signed W15TO10 = 0;
parameter signed W15TO11 = 0;
parameter signed W15TO12 = 0;
parameter signed W15TO13 = 0;
parameter signed W15TO14 = 0;
parameter signed W15TO15 = 0;
parameter signed W15TO16 = 0;
parameter signed W15TO17 = 0;
parameter signed W15TO18 = 0;
parameter signed W15TO19 = 0;
parameter signed W15TO20 = 0;
parameter signed W15TO21 = 0;
parameter signed W15TO22 = 0;
parameter signed W15TO23 = 0;
parameter signed W15TO24 = 0;
parameter signed W15TO25 = 0;
parameter signed W15TO26 = 0;
parameter signed W15TO27 = 0;
parameter signed W15TO28 = 0;
parameter signed W15TO29 = 0;
parameter signed W15TO30 = 0;
parameter signed W15TO31 = 0;
parameter signed W15TO32 = 0;
parameter signed W15TO33 = 0;
parameter signed W15TO34 = 0;
parameter signed W15TO35 = 0;
parameter signed W15TO36 = 0;
parameter signed W15TO37 = 0;
parameter signed W15TO38 = 0;
parameter signed W15TO39 = 0;
parameter signed W15TO40 = 0;
parameter signed W15TO41 = 0;
parameter signed W15TO42 = 0;
parameter signed W15TO43 = 0;
parameter signed W15TO44 = 0;
parameter signed W15TO45 = 0;
parameter signed W15TO46 = 0;
parameter signed W15TO47 = 0;
parameter signed W15TO48 = 0;
parameter signed W15TO49 = 0;
parameter signed W15TO50 = 0;
parameter signed W15TO51 = 0;
parameter signed W15TO52 = 0;
parameter signed W15TO53 = 0;
parameter signed W15TO54 = 0;
parameter signed W15TO55 = 0;
parameter signed W15TO56 = 0;
parameter signed W15TO57 = 0;
parameter signed W15TO58 = 0;
parameter signed W15TO59 = 0;
parameter signed W15TO60 = 0;
parameter signed W15TO61 = 0;
parameter signed W15TO62 = 0;
parameter signed W15TO63 = 0;
parameter signed W16TO0 = 0;
parameter signed W16TO1 = 0;
parameter signed W16TO2 = 0;
parameter signed W16TO3 = 0;
parameter signed W16TO4 = 0;
parameter signed W16TO5 = 0;
parameter signed W16TO6 = 0;
parameter signed W16TO7 = 0;
parameter signed W16TO8 = 0;
parameter signed W16TO9 = 0;
parameter signed W16TO10 = 0;
parameter signed W16TO11 = 0;
parameter signed W16TO12 = 0;
parameter signed W16TO13 = 0;
parameter signed W16TO14 = 0;
parameter signed W16TO15 = 0;
parameter signed W16TO16 = 0;
parameter signed W16TO17 = 0;
parameter signed W16TO18 = 0;
parameter signed W16TO19 = 0;
parameter signed W16TO20 = 0;
parameter signed W16TO21 = 0;
parameter signed W16TO22 = 0;
parameter signed W16TO23 = 0;
parameter signed W16TO24 = 0;
parameter signed W16TO25 = 0;
parameter signed W16TO26 = 0;
parameter signed W16TO27 = 0;
parameter signed W16TO28 = 0;
parameter signed W16TO29 = 0;
parameter signed W16TO30 = 0;
parameter signed W16TO31 = 0;
parameter signed W16TO32 = 0;
parameter signed W16TO33 = 0;
parameter signed W16TO34 = 0;
parameter signed W16TO35 = 0;
parameter signed W16TO36 = 0;
parameter signed W16TO37 = 0;
parameter signed W16TO38 = 0;
parameter signed W16TO39 = 0;
parameter signed W16TO40 = 0;
parameter signed W16TO41 = 0;
parameter signed W16TO42 = 0;
parameter signed W16TO43 = 0;
parameter signed W16TO44 = 0;
parameter signed W16TO45 = 0;
parameter signed W16TO46 = 0;
parameter signed W16TO47 = 0;
parameter signed W16TO48 = 0;
parameter signed W16TO49 = 0;
parameter signed W16TO50 = 0;
parameter signed W16TO51 = 0;
parameter signed W16TO52 = 0;
parameter signed W16TO53 = 0;
parameter signed W16TO54 = 0;
parameter signed W16TO55 = 0;
parameter signed W16TO56 = 0;
parameter signed W16TO57 = 0;
parameter signed W16TO58 = 0;
parameter signed W16TO59 = 0;
parameter signed W16TO60 = 0;
parameter signed W16TO61 = 0;
parameter signed W16TO62 = 0;
parameter signed W16TO63 = 0;
parameter signed W17TO0 = 0;
parameter signed W17TO1 = 0;
parameter signed W17TO2 = 0;
parameter signed W17TO3 = 0;
parameter signed W17TO4 = 0;
parameter signed W17TO5 = 0;
parameter signed W17TO6 = 0;
parameter signed W17TO7 = 0;
parameter signed W17TO8 = 0;
parameter signed W17TO9 = 0;
parameter signed W17TO10 = 0;
parameter signed W17TO11 = 0;
parameter signed W17TO12 = 0;
parameter signed W17TO13 = 0;
parameter signed W17TO14 = 0;
parameter signed W17TO15 = 0;
parameter signed W17TO16 = 0;
parameter signed W17TO17 = 0;
parameter signed W17TO18 = 0;
parameter signed W17TO19 = 0;
parameter signed W17TO20 = 0;
parameter signed W17TO21 = 0;
parameter signed W17TO22 = 0;
parameter signed W17TO23 = 0;
parameter signed W17TO24 = 0;
parameter signed W17TO25 = 0;
parameter signed W17TO26 = 0;
parameter signed W17TO27 = 0;
parameter signed W17TO28 = 0;
parameter signed W17TO29 = 0;
parameter signed W17TO30 = 0;
parameter signed W17TO31 = 0;
parameter signed W17TO32 = 0;
parameter signed W17TO33 = 0;
parameter signed W17TO34 = 0;
parameter signed W17TO35 = 0;
parameter signed W17TO36 = 0;
parameter signed W17TO37 = 0;
parameter signed W17TO38 = 0;
parameter signed W17TO39 = 0;
parameter signed W17TO40 = 0;
parameter signed W17TO41 = 0;
parameter signed W17TO42 = 0;
parameter signed W17TO43 = 0;
parameter signed W17TO44 = 0;
parameter signed W17TO45 = 0;
parameter signed W17TO46 = 0;
parameter signed W17TO47 = 0;
parameter signed W17TO48 = 0;
parameter signed W17TO49 = 0;
parameter signed W17TO50 = 0;
parameter signed W17TO51 = 0;
parameter signed W17TO52 = 0;
parameter signed W17TO53 = 0;
parameter signed W17TO54 = 0;
parameter signed W17TO55 = 0;
parameter signed W17TO56 = 0;
parameter signed W17TO57 = 0;
parameter signed W17TO58 = 0;
parameter signed W17TO59 = 0;
parameter signed W17TO60 = 0;
parameter signed W17TO61 = 0;
parameter signed W17TO62 = 0;
parameter signed W17TO63 = 0;
parameter signed W18TO0 = 0;
parameter signed W18TO1 = 0;
parameter signed W18TO2 = 0;
parameter signed W18TO3 = 0;
parameter signed W18TO4 = 0;
parameter signed W18TO5 = 0;
parameter signed W18TO6 = 0;
parameter signed W18TO7 = 0;
parameter signed W18TO8 = 0;
parameter signed W18TO9 = 0;
parameter signed W18TO10 = 0;
parameter signed W18TO11 = 0;
parameter signed W18TO12 = 0;
parameter signed W18TO13 = 0;
parameter signed W18TO14 = 0;
parameter signed W18TO15 = 0;
parameter signed W18TO16 = 0;
parameter signed W18TO17 = 0;
parameter signed W18TO18 = 0;
parameter signed W18TO19 = 0;
parameter signed W18TO20 = 0;
parameter signed W18TO21 = 0;
parameter signed W18TO22 = 0;
parameter signed W18TO23 = 0;
parameter signed W18TO24 = 0;
parameter signed W18TO25 = 0;
parameter signed W18TO26 = 0;
parameter signed W18TO27 = 0;
parameter signed W18TO28 = 0;
parameter signed W18TO29 = 0;
parameter signed W18TO30 = 0;
parameter signed W18TO31 = 0;
parameter signed W18TO32 = 0;
parameter signed W18TO33 = 0;
parameter signed W18TO34 = 0;
parameter signed W18TO35 = 0;
parameter signed W18TO36 = 0;
parameter signed W18TO37 = 0;
parameter signed W18TO38 = 0;
parameter signed W18TO39 = 0;
parameter signed W18TO40 = 0;
parameter signed W18TO41 = 0;
parameter signed W18TO42 = 0;
parameter signed W18TO43 = 0;
parameter signed W18TO44 = 0;
parameter signed W18TO45 = 0;
parameter signed W18TO46 = 0;
parameter signed W18TO47 = 0;
parameter signed W18TO48 = 0;
parameter signed W18TO49 = 0;
parameter signed W18TO50 = 0;
parameter signed W18TO51 = 0;
parameter signed W18TO52 = 0;
parameter signed W18TO53 = 0;
parameter signed W18TO54 = 0;
parameter signed W18TO55 = 0;
parameter signed W18TO56 = 0;
parameter signed W18TO57 = 0;
parameter signed W18TO58 = 0;
parameter signed W18TO59 = 0;
parameter signed W18TO60 = 0;
parameter signed W18TO61 = 0;
parameter signed W18TO62 = 0;
parameter signed W18TO63 = 0;
parameter signed W19TO0 = 0;
parameter signed W19TO1 = 0;
parameter signed W19TO2 = 0;
parameter signed W19TO3 = 0;
parameter signed W19TO4 = 0;
parameter signed W19TO5 = 0;
parameter signed W19TO6 = 0;
parameter signed W19TO7 = 0;
parameter signed W19TO8 = 0;
parameter signed W19TO9 = 0;
parameter signed W19TO10 = 0;
parameter signed W19TO11 = 0;
parameter signed W19TO12 = 0;
parameter signed W19TO13 = 0;
parameter signed W19TO14 = 0;
parameter signed W19TO15 = 0;
parameter signed W19TO16 = 0;
parameter signed W19TO17 = 0;
parameter signed W19TO18 = 0;
parameter signed W19TO19 = 0;
parameter signed W19TO20 = 0;
parameter signed W19TO21 = 0;
parameter signed W19TO22 = 0;
parameter signed W19TO23 = 0;
parameter signed W19TO24 = 0;
parameter signed W19TO25 = 0;
parameter signed W19TO26 = 0;
parameter signed W19TO27 = 0;
parameter signed W19TO28 = 0;
parameter signed W19TO29 = 0;
parameter signed W19TO30 = 0;
parameter signed W19TO31 = 0;
parameter signed W19TO32 = 0;
parameter signed W19TO33 = 0;
parameter signed W19TO34 = 0;
parameter signed W19TO35 = 0;
parameter signed W19TO36 = 0;
parameter signed W19TO37 = 0;
parameter signed W19TO38 = 0;
parameter signed W19TO39 = 0;
parameter signed W19TO40 = 0;
parameter signed W19TO41 = 0;
parameter signed W19TO42 = 0;
parameter signed W19TO43 = 0;
parameter signed W19TO44 = 0;
parameter signed W19TO45 = 0;
parameter signed W19TO46 = 0;
parameter signed W19TO47 = 0;
parameter signed W19TO48 = 0;
parameter signed W19TO49 = 0;
parameter signed W19TO50 = 0;
parameter signed W19TO51 = 0;
parameter signed W19TO52 = 0;
parameter signed W19TO53 = 0;
parameter signed W19TO54 = 0;
parameter signed W19TO55 = 0;
parameter signed W19TO56 = 0;
parameter signed W19TO57 = 0;
parameter signed W19TO58 = 0;
parameter signed W19TO59 = 0;
parameter signed W19TO60 = 0;
parameter signed W19TO61 = 0;
parameter signed W19TO62 = 0;
parameter signed W19TO63 = 0;
parameter signed W20TO0 = 0;
parameter signed W20TO1 = 0;
parameter signed W20TO2 = 0;
parameter signed W20TO3 = 0;
parameter signed W20TO4 = 0;
parameter signed W20TO5 = 0;
parameter signed W20TO6 = 0;
parameter signed W20TO7 = 0;
parameter signed W20TO8 = 0;
parameter signed W20TO9 = 0;
parameter signed W20TO10 = 0;
parameter signed W20TO11 = 0;
parameter signed W20TO12 = 0;
parameter signed W20TO13 = 0;
parameter signed W20TO14 = 0;
parameter signed W20TO15 = 0;
parameter signed W20TO16 = 0;
parameter signed W20TO17 = 0;
parameter signed W20TO18 = 0;
parameter signed W20TO19 = 0;
parameter signed W20TO20 = 0;
parameter signed W20TO21 = 0;
parameter signed W20TO22 = 0;
parameter signed W20TO23 = 0;
parameter signed W20TO24 = 0;
parameter signed W20TO25 = 0;
parameter signed W20TO26 = 0;
parameter signed W20TO27 = 0;
parameter signed W20TO28 = 0;
parameter signed W20TO29 = 0;
parameter signed W20TO30 = 0;
parameter signed W20TO31 = 0;
parameter signed W20TO32 = 0;
parameter signed W20TO33 = 0;
parameter signed W20TO34 = 0;
parameter signed W20TO35 = 0;
parameter signed W20TO36 = 0;
parameter signed W20TO37 = 0;
parameter signed W20TO38 = 0;
parameter signed W20TO39 = 0;
parameter signed W20TO40 = 0;
parameter signed W20TO41 = 0;
parameter signed W20TO42 = 0;
parameter signed W20TO43 = 0;
parameter signed W20TO44 = 0;
parameter signed W20TO45 = 0;
parameter signed W20TO46 = 0;
parameter signed W20TO47 = 0;
parameter signed W20TO48 = 0;
parameter signed W20TO49 = 0;
parameter signed W20TO50 = 0;
parameter signed W20TO51 = 0;
parameter signed W20TO52 = 0;
parameter signed W20TO53 = 0;
parameter signed W20TO54 = 0;
parameter signed W20TO55 = 0;
parameter signed W20TO56 = 0;
parameter signed W20TO57 = 0;
parameter signed W20TO58 = 0;
parameter signed W20TO59 = 0;
parameter signed W20TO60 = 0;
parameter signed W20TO61 = 0;
parameter signed W20TO62 = 0;
parameter signed W20TO63 = 0;
parameter signed W21TO0 = 0;
parameter signed W21TO1 = 0;
parameter signed W21TO2 = 0;
parameter signed W21TO3 = 0;
parameter signed W21TO4 = 0;
parameter signed W21TO5 = 0;
parameter signed W21TO6 = 0;
parameter signed W21TO7 = 0;
parameter signed W21TO8 = 0;
parameter signed W21TO9 = 0;
parameter signed W21TO10 = 0;
parameter signed W21TO11 = 0;
parameter signed W21TO12 = 0;
parameter signed W21TO13 = 0;
parameter signed W21TO14 = 0;
parameter signed W21TO15 = 0;
parameter signed W21TO16 = 0;
parameter signed W21TO17 = 0;
parameter signed W21TO18 = 0;
parameter signed W21TO19 = 0;
parameter signed W21TO20 = 0;
parameter signed W21TO21 = 0;
parameter signed W21TO22 = 0;
parameter signed W21TO23 = 0;
parameter signed W21TO24 = 0;
parameter signed W21TO25 = 0;
parameter signed W21TO26 = 0;
parameter signed W21TO27 = 0;
parameter signed W21TO28 = 0;
parameter signed W21TO29 = 0;
parameter signed W21TO30 = 0;
parameter signed W21TO31 = 0;
parameter signed W21TO32 = 0;
parameter signed W21TO33 = 0;
parameter signed W21TO34 = 0;
parameter signed W21TO35 = 0;
parameter signed W21TO36 = 0;
parameter signed W21TO37 = 0;
parameter signed W21TO38 = 0;
parameter signed W21TO39 = 0;
parameter signed W21TO40 = 0;
parameter signed W21TO41 = 0;
parameter signed W21TO42 = 0;
parameter signed W21TO43 = 0;
parameter signed W21TO44 = 0;
parameter signed W21TO45 = 0;
parameter signed W21TO46 = 0;
parameter signed W21TO47 = 0;
parameter signed W21TO48 = 0;
parameter signed W21TO49 = 0;
parameter signed W21TO50 = 0;
parameter signed W21TO51 = 0;
parameter signed W21TO52 = 0;
parameter signed W21TO53 = 0;
parameter signed W21TO54 = 0;
parameter signed W21TO55 = 0;
parameter signed W21TO56 = 0;
parameter signed W21TO57 = 0;
parameter signed W21TO58 = 0;
parameter signed W21TO59 = 0;
parameter signed W21TO60 = 0;
parameter signed W21TO61 = 0;
parameter signed W21TO62 = 0;
parameter signed W21TO63 = 0;
parameter signed W22TO0 = 0;
parameter signed W22TO1 = 0;
parameter signed W22TO2 = 0;
parameter signed W22TO3 = 0;
parameter signed W22TO4 = 0;
parameter signed W22TO5 = 0;
parameter signed W22TO6 = 0;
parameter signed W22TO7 = 0;
parameter signed W22TO8 = 0;
parameter signed W22TO9 = 0;
parameter signed W22TO10 = 0;
parameter signed W22TO11 = 0;
parameter signed W22TO12 = 0;
parameter signed W22TO13 = 0;
parameter signed W22TO14 = 0;
parameter signed W22TO15 = 0;
parameter signed W22TO16 = 0;
parameter signed W22TO17 = 0;
parameter signed W22TO18 = 0;
parameter signed W22TO19 = 0;
parameter signed W22TO20 = 0;
parameter signed W22TO21 = 0;
parameter signed W22TO22 = 0;
parameter signed W22TO23 = 0;
parameter signed W22TO24 = 0;
parameter signed W22TO25 = 0;
parameter signed W22TO26 = 0;
parameter signed W22TO27 = 0;
parameter signed W22TO28 = 0;
parameter signed W22TO29 = 0;
parameter signed W22TO30 = 0;
parameter signed W22TO31 = 0;
parameter signed W22TO32 = 0;
parameter signed W22TO33 = 0;
parameter signed W22TO34 = 0;
parameter signed W22TO35 = 0;
parameter signed W22TO36 = 0;
parameter signed W22TO37 = 0;
parameter signed W22TO38 = 0;
parameter signed W22TO39 = 0;
parameter signed W22TO40 = 0;
parameter signed W22TO41 = 0;
parameter signed W22TO42 = 0;
parameter signed W22TO43 = 0;
parameter signed W22TO44 = 0;
parameter signed W22TO45 = 0;
parameter signed W22TO46 = 0;
parameter signed W22TO47 = 0;
parameter signed W22TO48 = 0;
parameter signed W22TO49 = 0;
parameter signed W22TO50 = 0;
parameter signed W22TO51 = 0;
parameter signed W22TO52 = 0;
parameter signed W22TO53 = 0;
parameter signed W22TO54 = 0;
parameter signed W22TO55 = 0;
parameter signed W22TO56 = 0;
parameter signed W22TO57 = 0;
parameter signed W22TO58 = 0;
parameter signed W22TO59 = 0;
parameter signed W22TO60 = 0;
parameter signed W22TO61 = 0;
parameter signed W22TO62 = 0;
parameter signed W22TO63 = 0;
parameter signed W23TO0 = 0;
parameter signed W23TO1 = 0;
parameter signed W23TO2 = 0;
parameter signed W23TO3 = 0;
parameter signed W23TO4 = 0;
parameter signed W23TO5 = 0;
parameter signed W23TO6 = 0;
parameter signed W23TO7 = 0;
parameter signed W23TO8 = 0;
parameter signed W23TO9 = 0;
parameter signed W23TO10 = 0;
parameter signed W23TO11 = 0;
parameter signed W23TO12 = 0;
parameter signed W23TO13 = 0;
parameter signed W23TO14 = 0;
parameter signed W23TO15 = 0;
parameter signed W23TO16 = 0;
parameter signed W23TO17 = 0;
parameter signed W23TO18 = 0;
parameter signed W23TO19 = 0;
parameter signed W23TO20 = 0;
parameter signed W23TO21 = 0;
parameter signed W23TO22 = 0;
parameter signed W23TO23 = 0;
parameter signed W23TO24 = 0;
parameter signed W23TO25 = 0;
parameter signed W23TO26 = 0;
parameter signed W23TO27 = 0;
parameter signed W23TO28 = 0;
parameter signed W23TO29 = 0;
parameter signed W23TO30 = 0;
parameter signed W23TO31 = 0;
parameter signed W23TO32 = 0;
parameter signed W23TO33 = 0;
parameter signed W23TO34 = 0;
parameter signed W23TO35 = 0;
parameter signed W23TO36 = 0;
parameter signed W23TO37 = 0;
parameter signed W23TO38 = 0;
parameter signed W23TO39 = 0;
parameter signed W23TO40 = 0;
parameter signed W23TO41 = 0;
parameter signed W23TO42 = 0;
parameter signed W23TO43 = 0;
parameter signed W23TO44 = 0;
parameter signed W23TO45 = 0;
parameter signed W23TO46 = 0;
parameter signed W23TO47 = 0;
parameter signed W23TO48 = 0;
parameter signed W23TO49 = 0;
parameter signed W23TO50 = 0;
parameter signed W23TO51 = 0;
parameter signed W23TO52 = 0;
parameter signed W23TO53 = 0;
parameter signed W23TO54 = 0;
parameter signed W23TO55 = 0;
parameter signed W23TO56 = 0;
parameter signed W23TO57 = 0;
parameter signed W23TO58 = 0;
parameter signed W23TO59 = 0;
parameter signed W23TO60 = 0;
parameter signed W23TO61 = 0;
parameter signed W23TO62 = 0;
parameter signed W23TO63 = 0;
parameter signed W24TO0 = 0;
parameter signed W24TO1 = 0;
parameter signed W24TO2 = 0;
parameter signed W24TO3 = 0;
parameter signed W24TO4 = 0;
parameter signed W24TO5 = 0;
parameter signed W24TO6 = 0;
parameter signed W24TO7 = 0;
parameter signed W24TO8 = 0;
parameter signed W24TO9 = 0;
parameter signed W24TO10 = 0;
parameter signed W24TO11 = 0;
parameter signed W24TO12 = 0;
parameter signed W24TO13 = 0;
parameter signed W24TO14 = 0;
parameter signed W24TO15 = 0;
parameter signed W24TO16 = 0;
parameter signed W24TO17 = 0;
parameter signed W24TO18 = 0;
parameter signed W24TO19 = 0;
parameter signed W24TO20 = 0;
parameter signed W24TO21 = 0;
parameter signed W24TO22 = 0;
parameter signed W24TO23 = 0;
parameter signed W24TO24 = 0;
parameter signed W24TO25 = 0;
parameter signed W24TO26 = 0;
parameter signed W24TO27 = 0;
parameter signed W24TO28 = 0;
parameter signed W24TO29 = 0;
parameter signed W24TO30 = 0;
parameter signed W24TO31 = 0;
parameter signed W24TO32 = 0;
parameter signed W24TO33 = 0;
parameter signed W24TO34 = 0;
parameter signed W24TO35 = 0;
parameter signed W24TO36 = 0;
parameter signed W24TO37 = 0;
parameter signed W24TO38 = 0;
parameter signed W24TO39 = 0;
parameter signed W24TO40 = 0;
parameter signed W24TO41 = 0;
parameter signed W24TO42 = 0;
parameter signed W24TO43 = 0;
parameter signed W24TO44 = 0;
parameter signed W24TO45 = 0;
parameter signed W24TO46 = 0;
parameter signed W24TO47 = 0;
parameter signed W24TO48 = 0;
parameter signed W24TO49 = 0;
parameter signed W24TO50 = 0;
parameter signed W24TO51 = 0;
parameter signed W24TO52 = 0;
parameter signed W24TO53 = 0;
parameter signed W24TO54 = 0;
parameter signed W24TO55 = 0;
parameter signed W24TO56 = 0;
parameter signed W24TO57 = 0;
parameter signed W24TO58 = 0;
parameter signed W24TO59 = 0;
parameter signed W24TO60 = 0;
parameter signed W24TO61 = 0;
parameter signed W24TO62 = 0;
parameter signed W24TO63 = 0;
parameter signed W25TO0 = 0;
parameter signed W25TO1 = 0;
parameter signed W25TO2 = 0;
parameter signed W25TO3 = 0;
parameter signed W25TO4 = 0;
parameter signed W25TO5 = 0;
parameter signed W25TO6 = 0;
parameter signed W25TO7 = 0;
parameter signed W25TO8 = 0;
parameter signed W25TO9 = 0;
parameter signed W25TO10 = 0;
parameter signed W25TO11 = 0;
parameter signed W25TO12 = 0;
parameter signed W25TO13 = 0;
parameter signed W25TO14 = 0;
parameter signed W25TO15 = 0;
parameter signed W25TO16 = 0;
parameter signed W25TO17 = 0;
parameter signed W25TO18 = 0;
parameter signed W25TO19 = 0;
parameter signed W25TO20 = 0;
parameter signed W25TO21 = 0;
parameter signed W25TO22 = 0;
parameter signed W25TO23 = 0;
parameter signed W25TO24 = 0;
parameter signed W25TO25 = 0;
parameter signed W25TO26 = 0;
parameter signed W25TO27 = 0;
parameter signed W25TO28 = 0;
parameter signed W25TO29 = 0;
parameter signed W25TO30 = 0;
parameter signed W25TO31 = 0;
parameter signed W25TO32 = 0;
parameter signed W25TO33 = 0;
parameter signed W25TO34 = 0;
parameter signed W25TO35 = 0;
parameter signed W25TO36 = 0;
parameter signed W25TO37 = 0;
parameter signed W25TO38 = 0;
parameter signed W25TO39 = 0;
parameter signed W25TO40 = 0;
parameter signed W25TO41 = 0;
parameter signed W25TO42 = 0;
parameter signed W25TO43 = 0;
parameter signed W25TO44 = 0;
parameter signed W25TO45 = 0;
parameter signed W25TO46 = 0;
parameter signed W25TO47 = 0;
parameter signed W25TO48 = 0;
parameter signed W25TO49 = 0;
parameter signed W25TO50 = 0;
parameter signed W25TO51 = 0;
parameter signed W25TO52 = 0;
parameter signed W25TO53 = 0;
parameter signed W25TO54 = 0;
parameter signed W25TO55 = 0;
parameter signed W25TO56 = 0;
parameter signed W25TO57 = 0;
parameter signed W25TO58 = 0;
parameter signed W25TO59 = 0;
parameter signed W25TO60 = 0;
parameter signed W25TO61 = 0;
parameter signed W25TO62 = 0;
parameter signed W25TO63 = 0;
parameter signed W26TO0 = 0;
parameter signed W26TO1 = 0;
parameter signed W26TO2 = 0;
parameter signed W26TO3 = 0;
parameter signed W26TO4 = 0;
parameter signed W26TO5 = 0;
parameter signed W26TO6 = 0;
parameter signed W26TO7 = 0;
parameter signed W26TO8 = 0;
parameter signed W26TO9 = 0;
parameter signed W26TO10 = 0;
parameter signed W26TO11 = 0;
parameter signed W26TO12 = 0;
parameter signed W26TO13 = 0;
parameter signed W26TO14 = 0;
parameter signed W26TO15 = 0;
parameter signed W26TO16 = 0;
parameter signed W26TO17 = 0;
parameter signed W26TO18 = 0;
parameter signed W26TO19 = 0;
parameter signed W26TO20 = 0;
parameter signed W26TO21 = 0;
parameter signed W26TO22 = 0;
parameter signed W26TO23 = 0;
parameter signed W26TO24 = 0;
parameter signed W26TO25 = 0;
parameter signed W26TO26 = 0;
parameter signed W26TO27 = 0;
parameter signed W26TO28 = 0;
parameter signed W26TO29 = 0;
parameter signed W26TO30 = 0;
parameter signed W26TO31 = 0;
parameter signed W26TO32 = 0;
parameter signed W26TO33 = 0;
parameter signed W26TO34 = 0;
parameter signed W26TO35 = 0;
parameter signed W26TO36 = 0;
parameter signed W26TO37 = 0;
parameter signed W26TO38 = 0;
parameter signed W26TO39 = 0;
parameter signed W26TO40 = 0;
parameter signed W26TO41 = 0;
parameter signed W26TO42 = 0;
parameter signed W26TO43 = 0;
parameter signed W26TO44 = 0;
parameter signed W26TO45 = 0;
parameter signed W26TO46 = 0;
parameter signed W26TO47 = 0;
parameter signed W26TO48 = 0;
parameter signed W26TO49 = 0;
parameter signed W26TO50 = 0;
parameter signed W26TO51 = 0;
parameter signed W26TO52 = 0;
parameter signed W26TO53 = 0;
parameter signed W26TO54 = 0;
parameter signed W26TO55 = 0;
parameter signed W26TO56 = 0;
parameter signed W26TO57 = 0;
parameter signed W26TO58 = 0;
parameter signed W26TO59 = 0;
parameter signed W26TO60 = 0;
parameter signed W26TO61 = 0;
parameter signed W26TO62 = 0;
parameter signed W26TO63 = 0;
parameter signed W27TO0 = 0;
parameter signed W27TO1 = 0;
parameter signed W27TO2 = 0;
parameter signed W27TO3 = 0;
parameter signed W27TO4 = 0;
parameter signed W27TO5 = 0;
parameter signed W27TO6 = 0;
parameter signed W27TO7 = 0;
parameter signed W27TO8 = 0;
parameter signed W27TO9 = 0;
parameter signed W27TO10 = 0;
parameter signed W27TO11 = 0;
parameter signed W27TO12 = 0;
parameter signed W27TO13 = 0;
parameter signed W27TO14 = 0;
parameter signed W27TO15 = 0;
parameter signed W27TO16 = 0;
parameter signed W27TO17 = 0;
parameter signed W27TO18 = 0;
parameter signed W27TO19 = 0;
parameter signed W27TO20 = 0;
parameter signed W27TO21 = 0;
parameter signed W27TO22 = 0;
parameter signed W27TO23 = 0;
parameter signed W27TO24 = 0;
parameter signed W27TO25 = 0;
parameter signed W27TO26 = 0;
parameter signed W27TO27 = 0;
parameter signed W27TO28 = 0;
parameter signed W27TO29 = 0;
parameter signed W27TO30 = 0;
parameter signed W27TO31 = 0;
parameter signed W27TO32 = 0;
parameter signed W27TO33 = 0;
parameter signed W27TO34 = 0;
parameter signed W27TO35 = 0;
parameter signed W27TO36 = 0;
parameter signed W27TO37 = 0;
parameter signed W27TO38 = 0;
parameter signed W27TO39 = 0;
parameter signed W27TO40 = 0;
parameter signed W27TO41 = 0;
parameter signed W27TO42 = 0;
parameter signed W27TO43 = 0;
parameter signed W27TO44 = 0;
parameter signed W27TO45 = 0;
parameter signed W27TO46 = 0;
parameter signed W27TO47 = 0;
parameter signed W27TO48 = 0;
parameter signed W27TO49 = 0;
parameter signed W27TO50 = 0;
parameter signed W27TO51 = 0;
parameter signed W27TO52 = 0;
parameter signed W27TO53 = 0;
parameter signed W27TO54 = 0;
parameter signed W27TO55 = 0;
parameter signed W27TO56 = 0;
parameter signed W27TO57 = 0;
parameter signed W27TO58 = 0;
parameter signed W27TO59 = 0;
parameter signed W27TO60 = 0;
parameter signed W27TO61 = 0;
parameter signed W27TO62 = 0;
parameter signed W27TO63 = 0;
parameter signed W28TO0 = 0;
parameter signed W28TO1 = 0;
parameter signed W28TO2 = 0;
parameter signed W28TO3 = 0;
parameter signed W28TO4 = 0;
parameter signed W28TO5 = 0;
parameter signed W28TO6 = 0;
parameter signed W28TO7 = 0;
parameter signed W28TO8 = 0;
parameter signed W28TO9 = 0;
parameter signed W28TO10 = 0;
parameter signed W28TO11 = 0;
parameter signed W28TO12 = 0;
parameter signed W28TO13 = 0;
parameter signed W28TO14 = 0;
parameter signed W28TO15 = 0;
parameter signed W28TO16 = 0;
parameter signed W28TO17 = 0;
parameter signed W28TO18 = 0;
parameter signed W28TO19 = 0;
parameter signed W28TO20 = 0;
parameter signed W28TO21 = 0;
parameter signed W28TO22 = 0;
parameter signed W28TO23 = 0;
parameter signed W28TO24 = 0;
parameter signed W28TO25 = 0;
parameter signed W28TO26 = 0;
parameter signed W28TO27 = 0;
parameter signed W28TO28 = 0;
parameter signed W28TO29 = 0;
parameter signed W28TO30 = 0;
parameter signed W28TO31 = 0;
parameter signed W28TO32 = 0;
parameter signed W28TO33 = 0;
parameter signed W28TO34 = 0;
parameter signed W28TO35 = 0;
parameter signed W28TO36 = 0;
parameter signed W28TO37 = 0;
parameter signed W28TO38 = 0;
parameter signed W28TO39 = 0;
parameter signed W28TO40 = 0;
parameter signed W28TO41 = 0;
parameter signed W28TO42 = 0;
parameter signed W28TO43 = 0;
parameter signed W28TO44 = 0;
parameter signed W28TO45 = 0;
parameter signed W28TO46 = 0;
parameter signed W28TO47 = 0;
parameter signed W28TO48 = 0;
parameter signed W28TO49 = 0;
parameter signed W28TO50 = 0;
parameter signed W28TO51 = 0;
parameter signed W28TO52 = 0;
parameter signed W28TO53 = 0;
parameter signed W28TO54 = 0;
parameter signed W28TO55 = 0;
parameter signed W28TO56 = 0;
parameter signed W28TO57 = 0;
parameter signed W28TO58 = 0;
parameter signed W28TO59 = 0;
parameter signed W28TO60 = 0;
parameter signed W28TO61 = 0;
parameter signed W28TO62 = 0;
parameter signed W28TO63 = 0;
parameter signed W29TO0 = 0;
parameter signed W29TO1 = 0;
parameter signed W29TO2 = 0;
parameter signed W29TO3 = 0;
parameter signed W29TO4 = 0;
parameter signed W29TO5 = 0;
parameter signed W29TO6 = 0;
parameter signed W29TO7 = 0;
parameter signed W29TO8 = 0;
parameter signed W29TO9 = 0;
parameter signed W29TO10 = 0;
parameter signed W29TO11 = 0;
parameter signed W29TO12 = 0;
parameter signed W29TO13 = 0;
parameter signed W29TO14 = 0;
parameter signed W29TO15 = 0;
parameter signed W29TO16 = 0;
parameter signed W29TO17 = 0;
parameter signed W29TO18 = 0;
parameter signed W29TO19 = 0;
parameter signed W29TO20 = 0;
parameter signed W29TO21 = 0;
parameter signed W29TO22 = 0;
parameter signed W29TO23 = 0;
parameter signed W29TO24 = 0;
parameter signed W29TO25 = 0;
parameter signed W29TO26 = 0;
parameter signed W29TO27 = 0;
parameter signed W29TO28 = 0;
parameter signed W29TO29 = 0;
parameter signed W29TO30 = 0;
parameter signed W29TO31 = 0;
parameter signed W29TO32 = 0;
parameter signed W29TO33 = 0;
parameter signed W29TO34 = 0;
parameter signed W29TO35 = 0;
parameter signed W29TO36 = 0;
parameter signed W29TO37 = 0;
parameter signed W29TO38 = 0;
parameter signed W29TO39 = 0;
parameter signed W29TO40 = 0;
parameter signed W29TO41 = 0;
parameter signed W29TO42 = 0;
parameter signed W29TO43 = 0;
parameter signed W29TO44 = 0;
parameter signed W29TO45 = 0;
parameter signed W29TO46 = 0;
parameter signed W29TO47 = 0;
parameter signed W29TO48 = 0;
parameter signed W29TO49 = 0;
parameter signed W29TO50 = 0;
parameter signed W29TO51 = 0;
parameter signed W29TO52 = 0;
parameter signed W29TO53 = 0;
parameter signed W29TO54 = 0;
parameter signed W29TO55 = 0;
parameter signed W29TO56 = 0;
parameter signed W29TO57 = 0;
parameter signed W29TO58 = 0;
parameter signed W29TO59 = 0;
parameter signed W29TO60 = 0;
parameter signed W29TO61 = 0;
parameter signed W29TO62 = 0;
parameter signed W29TO63 = 0;
parameter signed W30TO0 = 0;
parameter signed W30TO1 = 0;
parameter signed W30TO2 = 0;
parameter signed W30TO3 = 0;
parameter signed W30TO4 = 0;
parameter signed W30TO5 = 0;
parameter signed W30TO6 = 0;
parameter signed W30TO7 = 0;
parameter signed W30TO8 = 0;
parameter signed W30TO9 = 0;
parameter signed W30TO10 = 0;
parameter signed W30TO11 = 0;
parameter signed W30TO12 = 0;
parameter signed W30TO13 = 0;
parameter signed W30TO14 = 0;
parameter signed W30TO15 = 0;
parameter signed W30TO16 = 0;
parameter signed W30TO17 = 0;
parameter signed W30TO18 = 0;
parameter signed W30TO19 = 0;
parameter signed W30TO20 = 0;
parameter signed W30TO21 = 0;
parameter signed W30TO22 = 0;
parameter signed W30TO23 = 0;
parameter signed W30TO24 = 0;
parameter signed W30TO25 = 0;
parameter signed W30TO26 = 0;
parameter signed W30TO27 = 0;
parameter signed W30TO28 = 0;
parameter signed W30TO29 = 0;
parameter signed W30TO30 = 0;
parameter signed W30TO31 = 0;
parameter signed W30TO32 = 0;
parameter signed W30TO33 = 0;
parameter signed W30TO34 = 0;
parameter signed W30TO35 = 0;
parameter signed W30TO36 = 0;
parameter signed W30TO37 = 0;
parameter signed W30TO38 = 0;
parameter signed W30TO39 = 0;
parameter signed W30TO40 = 0;
parameter signed W30TO41 = 0;
parameter signed W30TO42 = 0;
parameter signed W30TO43 = 0;
parameter signed W30TO44 = 0;
parameter signed W30TO45 = 0;
parameter signed W30TO46 = 0;
parameter signed W30TO47 = 0;
parameter signed W30TO48 = 0;
parameter signed W30TO49 = 0;
parameter signed W30TO50 = 0;
parameter signed W30TO51 = 0;
parameter signed W30TO52 = 0;
parameter signed W30TO53 = 0;
parameter signed W30TO54 = 0;
parameter signed W30TO55 = 0;
parameter signed W30TO56 = 0;
parameter signed W30TO57 = 0;
parameter signed W30TO58 = 0;
parameter signed W30TO59 = 0;
parameter signed W30TO60 = 0;
parameter signed W30TO61 = 0;
parameter signed W30TO62 = 0;
parameter signed W30TO63 = 0;
parameter signed W31TO0 = 0;
parameter signed W31TO1 = 0;
parameter signed W31TO2 = 0;
parameter signed W31TO3 = 0;
parameter signed W31TO4 = 0;
parameter signed W31TO5 = 0;
parameter signed W31TO6 = 0;
parameter signed W31TO7 = 0;
parameter signed W31TO8 = 0;
parameter signed W31TO9 = 0;
parameter signed W31TO10 = 0;
parameter signed W31TO11 = 0;
parameter signed W31TO12 = 0;
parameter signed W31TO13 = 0;
parameter signed W31TO14 = 0;
parameter signed W31TO15 = 0;
parameter signed W31TO16 = 0;
parameter signed W31TO17 = 0;
parameter signed W31TO18 = 0;
parameter signed W31TO19 = 0;
parameter signed W31TO20 = 0;
parameter signed W31TO21 = 0;
parameter signed W31TO22 = 0;
parameter signed W31TO23 = 0;
parameter signed W31TO24 = 0;
parameter signed W31TO25 = 0;
parameter signed W31TO26 = 0;
parameter signed W31TO27 = 0;
parameter signed W31TO28 = 0;
parameter signed W31TO29 = 0;
parameter signed W31TO30 = 0;
parameter signed W31TO31 = 0;
parameter signed W31TO32 = 0;
parameter signed W31TO33 = 0;
parameter signed W31TO34 = 0;
parameter signed W31TO35 = 0;
parameter signed W31TO36 = 0;
parameter signed W31TO37 = 0;
parameter signed W31TO38 = 0;
parameter signed W31TO39 = 0;
parameter signed W31TO40 = 0;
parameter signed W31TO41 = 0;
parameter signed W31TO42 = 0;
parameter signed W31TO43 = 0;
parameter signed W31TO44 = 0;
parameter signed W31TO45 = 0;
parameter signed W31TO46 = 0;
parameter signed W31TO47 = 0;
parameter signed W31TO48 = 0;
parameter signed W31TO49 = 0;
parameter signed W31TO50 = 0;
parameter signed W31TO51 = 0;
parameter signed W31TO52 = 0;
parameter signed W31TO53 = 0;
parameter signed W31TO54 = 0;
parameter signed W31TO55 = 0;
parameter signed W31TO56 = 0;
parameter signed W31TO57 = 0;
parameter signed W31TO58 = 0;
parameter signed W31TO59 = 0;
parameter signed W31TO60 = 0;
parameter signed W31TO61 = 0;
parameter signed W31TO62 = 0;
parameter signed W31TO63 = 0;
parameter signed W32TO0 = 0;
parameter signed W32TO1 = 0;
parameter signed W32TO2 = 0;
parameter signed W32TO3 = 0;
parameter signed W32TO4 = 0;
parameter signed W32TO5 = 0;
parameter signed W32TO6 = 0;
parameter signed W32TO7 = 0;
parameter signed W32TO8 = 0;
parameter signed W32TO9 = 0;
parameter signed W32TO10 = 0;
parameter signed W32TO11 = 0;
parameter signed W32TO12 = 0;
parameter signed W32TO13 = 0;
parameter signed W32TO14 = 0;
parameter signed W32TO15 = 0;
parameter signed W32TO16 = 0;
parameter signed W32TO17 = 0;
parameter signed W32TO18 = 0;
parameter signed W32TO19 = 0;
parameter signed W32TO20 = 0;
parameter signed W32TO21 = 0;
parameter signed W32TO22 = 0;
parameter signed W32TO23 = 0;
parameter signed W32TO24 = 0;
parameter signed W32TO25 = 0;
parameter signed W32TO26 = 0;
parameter signed W32TO27 = 0;
parameter signed W32TO28 = 0;
parameter signed W32TO29 = 0;
parameter signed W32TO30 = 0;
parameter signed W32TO31 = 0;
parameter signed W32TO32 = 0;
parameter signed W32TO33 = 0;
parameter signed W32TO34 = 0;
parameter signed W32TO35 = 0;
parameter signed W32TO36 = 0;
parameter signed W32TO37 = 0;
parameter signed W32TO38 = 0;
parameter signed W32TO39 = 0;
parameter signed W32TO40 = 0;
parameter signed W32TO41 = 0;
parameter signed W32TO42 = 0;
parameter signed W32TO43 = 0;
parameter signed W32TO44 = 0;
parameter signed W32TO45 = 0;
parameter signed W32TO46 = 0;
parameter signed W32TO47 = 0;
parameter signed W32TO48 = 0;
parameter signed W32TO49 = 0;
parameter signed W32TO50 = 0;
parameter signed W32TO51 = 0;
parameter signed W32TO52 = 0;
parameter signed W32TO53 = 0;
parameter signed W32TO54 = 0;
parameter signed W32TO55 = 0;
parameter signed W32TO56 = 0;
parameter signed W32TO57 = 0;
parameter signed W32TO58 = 0;
parameter signed W32TO59 = 0;
parameter signed W32TO60 = 0;
parameter signed W32TO61 = 0;
parameter signed W32TO62 = 0;
parameter signed W32TO63 = 0;
parameter signed W33TO0 = 0;
parameter signed W33TO1 = 0;
parameter signed W33TO2 = 0;
parameter signed W33TO3 = 0;
parameter signed W33TO4 = 0;
parameter signed W33TO5 = 0;
parameter signed W33TO6 = 0;
parameter signed W33TO7 = 0;
parameter signed W33TO8 = 0;
parameter signed W33TO9 = 0;
parameter signed W33TO10 = 0;
parameter signed W33TO11 = 0;
parameter signed W33TO12 = 0;
parameter signed W33TO13 = 0;
parameter signed W33TO14 = 0;
parameter signed W33TO15 = 0;
parameter signed W33TO16 = 0;
parameter signed W33TO17 = 0;
parameter signed W33TO18 = 0;
parameter signed W33TO19 = 0;
parameter signed W33TO20 = 0;
parameter signed W33TO21 = 0;
parameter signed W33TO22 = 0;
parameter signed W33TO23 = 0;
parameter signed W33TO24 = 0;
parameter signed W33TO25 = 0;
parameter signed W33TO26 = 0;
parameter signed W33TO27 = 0;
parameter signed W33TO28 = 0;
parameter signed W33TO29 = 0;
parameter signed W33TO30 = 0;
parameter signed W33TO31 = 0;
parameter signed W33TO32 = 0;
parameter signed W33TO33 = 0;
parameter signed W33TO34 = 0;
parameter signed W33TO35 = 0;
parameter signed W33TO36 = 0;
parameter signed W33TO37 = 0;
parameter signed W33TO38 = 0;
parameter signed W33TO39 = 0;
parameter signed W33TO40 = 0;
parameter signed W33TO41 = 0;
parameter signed W33TO42 = 0;
parameter signed W33TO43 = 0;
parameter signed W33TO44 = 0;
parameter signed W33TO45 = 0;
parameter signed W33TO46 = 0;
parameter signed W33TO47 = 0;
parameter signed W33TO48 = 0;
parameter signed W33TO49 = 0;
parameter signed W33TO50 = 0;
parameter signed W33TO51 = 0;
parameter signed W33TO52 = 0;
parameter signed W33TO53 = 0;
parameter signed W33TO54 = 0;
parameter signed W33TO55 = 0;
parameter signed W33TO56 = 0;
parameter signed W33TO57 = 0;
parameter signed W33TO58 = 0;
parameter signed W33TO59 = 0;
parameter signed W33TO60 = 0;
parameter signed W33TO61 = 0;
parameter signed W33TO62 = 0;
parameter signed W33TO63 = 0;
parameter signed W34TO0 = 0;
parameter signed W34TO1 = 0;
parameter signed W34TO2 = 0;
parameter signed W34TO3 = 0;
parameter signed W34TO4 = 0;
parameter signed W34TO5 = 0;
parameter signed W34TO6 = 0;
parameter signed W34TO7 = 0;
parameter signed W34TO8 = 0;
parameter signed W34TO9 = 0;
parameter signed W34TO10 = 0;
parameter signed W34TO11 = 0;
parameter signed W34TO12 = 0;
parameter signed W34TO13 = 0;
parameter signed W34TO14 = 0;
parameter signed W34TO15 = 0;
parameter signed W34TO16 = 0;
parameter signed W34TO17 = 0;
parameter signed W34TO18 = 0;
parameter signed W34TO19 = 0;
parameter signed W34TO20 = 0;
parameter signed W34TO21 = 0;
parameter signed W34TO22 = 0;
parameter signed W34TO23 = 0;
parameter signed W34TO24 = 0;
parameter signed W34TO25 = 0;
parameter signed W34TO26 = 0;
parameter signed W34TO27 = 0;
parameter signed W34TO28 = 0;
parameter signed W34TO29 = 0;
parameter signed W34TO30 = 0;
parameter signed W34TO31 = 0;
parameter signed W34TO32 = 0;
parameter signed W34TO33 = 0;
parameter signed W34TO34 = 0;
parameter signed W34TO35 = 0;
parameter signed W34TO36 = 0;
parameter signed W34TO37 = 0;
parameter signed W34TO38 = 0;
parameter signed W34TO39 = 0;
parameter signed W34TO40 = 0;
parameter signed W34TO41 = 0;
parameter signed W34TO42 = 0;
parameter signed W34TO43 = 0;
parameter signed W34TO44 = 0;
parameter signed W34TO45 = 0;
parameter signed W34TO46 = 0;
parameter signed W34TO47 = 0;
parameter signed W34TO48 = 0;
parameter signed W34TO49 = 0;
parameter signed W34TO50 = 0;
parameter signed W34TO51 = 0;
parameter signed W34TO52 = 0;
parameter signed W34TO53 = 0;
parameter signed W34TO54 = 0;
parameter signed W34TO55 = 0;
parameter signed W34TO56 = 0;
parameter signed W34TO57 = 0;
parameter signed W34TO58 = 0;
parameter signed W34TO59 = 0;
parameter signed W34TO60 = 0;
parameter signed W34TO61 = 0;
parameter signed W34TO62 = 0;
parameter signed W34TO63 = 0;
parameter signed W35TO0 = 0;
parameter signed W35TO1 = 0;
parameter signed W35TO2 = 0;
parameter signed W35TO3 = 0;
parameter signed W35TO4 = 0;
parameter signed W35TO5 = 0;
parameter signed W35TO6 = 0;
parameter signed W35TO7 = 0;
parameter signed W35TO8 = 0;
parameter signed W35TO9 = 0;
parameter signed W35TO10 = 0;
parameter signed W35TO11 = 0;
parameter signed W35TO12 = 0;
parameter signed W35TO13 = 0;
parameter signed W35TO14 = 0;
parameter signed W35TO15 = 0;
parameter signed W35TO16 = 0;
parameter signed W35TO17 = 0;
parameter signed W35TO18 = 0;
parameter signed W35TO19 = 0;
parameter signed W35TO20 = 0;
parameter signed W35TO21 = 0;
parameter signed W35TO22 = 0;
parameter signed W35TO23 = 0;
parameter signed W35TO24 = 0;
parameter signed W35TO25 = 0;
parameter signed W35TO26 = 0;
parameter signed W35TO27 = 0;
parameter signed W35TO28 = 0;
parameter signed W35TO29 = 0;
parameter signed W35TO30 = 0;
parameter signed W35TO31 = 0;
parameter signed W35TO32 = 0;
parameter signed W35TO33 = 0;
parameter signed W35TO34 = 0;
parameter signed W35TO35 = 0;
parameter signed W35TO36 = 0;
parameter signed W35TO37 = 0;
parameter signed W35TO38 = 0;
parameter signed W35TO39 = 0;
parameter signed W35TO40 = 0;
parameter signed W35TO41 = 0;
parameter signed W35TO42 = 0;
parameter signed W35TO43 = 0;
parameter signed W35TO44 = 0;
parameter signed W35TO45 = 0;
parameter signed W35TO46 = 0;
parameter signed W35TO47 = 0;
parameter signed W35TO48 = 0;
parameter signed W35TO49 = 0;
parameter signed W35TO50 = 0;
parameter signed W35TO51 = 0;
parameter signed W35TO52 = 0;
parameter signed W35TO53 = 0;
parameter signed W35TO54 = 0;
parameter signed W35TO55 = 0;
parameter signed W35TO56 = 0;
parameter signed W35TO57 = 0;
parameter signed W35TO58 = 0;
parameter signed W35TO59 = 0;
parameter signed W35TO60 = 0;
parameter signed W35TO61 = 0;
parameter signed W35TO62 = 0;
parameter signed W35TO63 = 0;
parameter signed W36TO0 = 0;
parameter signed W36TO1 = 0;
parameter signed W36TO2 = 0;
parameter signed W36TO3 = 0;
parameter signed W36TO4 = 0;
parameter signed W36TO5 = 0;
parameter signed W36TO6 = 0;
parameter signed W36TO7 = 0;
parameter signed W36TO8 = 0;
parameter signed W36TO9 = 0;
parameter signed W36TO10 = 0;
parameter signed W36TO11 = 0;
parameter signed W36TO12 = 0;
parameter signed W36TO13 = 0;
parameter signed W36TO14 = 0;
parameter signed W36TO15 = 0;
parameter signed W36TO16 = 0;
parameter signed W36TO17 = 0;
parameter signed W36TO18 = 0;
parameter signed W36TO19 = 0;
parameter signed W36TO20 = 0;
parameter signed W36TO21 = 0;
parameter signed W36TO22 = 0;
parameter signed W36TO23 = 0;
parameter signed W36TO24 = 0;
parameter signed W36TO25 = 0;
parameter signed W36TO26 = 0;
parameter signed W36TO27 = 0;
parameter signed W36TO28 = 0;
parameter signed W36TO29 = 0;
parameter signed W36TO30 = 0;
parameter signed W36TO31 = 0;
parameter signed W36TO32 = 0;
parameter signed W36TO33 = 0;
parameter signed W36TO34 = 0;
parameter signed W36TO35 = 0;
parameter signed W36TO36 = 0;
parameter signed W36TO37 = 0;
parameter signed W36TO38 = 0;
parameter signed W36TO39 = 0;
parameter signed W36TO40 = 0;
parameter signed W36TO41 = 0;
parameter signed W36TO42 = 0;
parameter signed W36TO43 = 0;
parameter signed W36TO44 = 0;
parameter signed W36TO45 = 0;
parameter signed W36TO46 = 0;
parameter signed W36TO47 = 0;
parameter signed W36TO48 = 0;
parameter signed W36TO49 = 0;
parameter signed W36TO50 = 0;
parameter signed W36TO51 = 0;
parameter signed W36TO52 = 0;
parameter signed W36TO53 = 0;
parameter signed W36TO54 = 0;
parameter signed W36TO55 = 0;
parameter signed W36TO56 = 0;
parameter signed W36TO57 = 0;
parameter signed W36TO58 = 0;
parameter signed W36TO59 = 0;
parameter signed W36TO60 = 0;
parameter signed W36TO61 = 0;
parameter signed W36TO62 = 0;
parameter signed W36TO63 = 0;
parameter signed W37TO0 = 0;
parameter signed W37TO1 = 0;
parameter signed W37TO2 = 0;
parameter signed W37TO3 = 0;
parameter signed W37TO4 = 0;
parameter signed W37TO5 = 0;
parameter signed W37TO6 = 0;
parameter signed W37TO7 = 0;
parameter signed W37TO8 = 0;
parameter signed W37TO9 = 0;
parameter signed W37TO10 = 0;
parameter signed W37TO11 = 0;
parameter signed W37TO12 = 0;
parameter signed W37TO13 = 0;
parameter signed W37TO14 = 0;
parameter signed W37TO15 = 0;
parameter signed W37TO16 = 0;
parameter signed W37TO17 = 0;
parameter signed W37TO18 = 0;
parameter signed W37TO19 = 0;
parameter signed W37TO20 = 0;
parameter signed W37TO21 = 0;
parameter signed W37TO22 = 0;
parameter signed W37TO23 = 0;
parameter signed W37TO24 = 0;
parameter signed W37TO25 = 0;
parameter signed W37TO26 = 0;
parameter signed W37TO27 = 0;
parameter signed W37TO28 = 0;
parameter signed W37TO29 = 0;
parameter signed W37TO30 = 0;
parameter signed W37TO31 = 0;
parameter signed W37TO32 = 0;
parameter signed W37TO33 = 0;
parameter signed W37TO34 = 0;
parameter signed W37TO35 = 0;
parameter signed W37TO36 = 0;
parameter signed W37TO37 = 0;
parameter signed W37TO38 = 0;
parameter signed W37TO39 = 0;
parameter signed W37TO40 = 0;
parameter signed W37TO41 = 0;
parameter signed W37TO42 = 0;
parameter signed W37TO43 = 0;
parameter signed W37TO44 = 0;
parameter signed W37TO45 = 0;
parameter signed W37TO46 = 0;
parameter signed W37TO47 = 0;
parameter signed W37TO48 = 0;
parameter signed W37TO49 = 0;
parameter signed W37TO50 = 0;
parameter signed W37TO51 = 0;
parameter signed W37TO52 = 0;
parameter signed W37TO53 = 0;
parameter signed W37TO54 = 0;
parameter signed W37TO55 = 0;
parameter signed W37TO56 = 0;
parameter signed W37TO57 = 0;
parameter signed W37TO58 = 0;
parameter signed W37TO59 = 0;
parameter signed W37TO60 = 0;
parameter signed W37TO61 = 0;
parameter signed W37TO62 = 0;
parameter signed W37TO63 = 0;
parameter signed W38TO0 = 0;
parameter signed W38TO1 = 0;
parameter signed W38TO2 = 0;
parameter signed W38TO3 = 0;
parameter signed W38TO4 = 0;
parameter signed W38TO5 = 0;
parameter signed W38TO6 = 0;
parameter signed W38TO7 = 0;
parameter signed W38TO8 = 0;
parameter signed W38TO9 = 0;
parameter signed W38TO10 = 0;
parameter signed W38TO11 = 0;
parameter signed W38TO12 = 0;
parameter signed W38TO13 = 0;
parameter signed W38TO14 = 0;
parameter signed W38TO15 = 0;
parameter signed W38TO16 = 0;
parameter signed W38TO17 = 0;
parameter signed W38TO18 = 0;
parameter signed W38TO19 = 0;
parameter signed W38TO20 = 0;
parameter signed W38TO21 = 0;
parameter signed W38TO22 = 0;
parameter signed W38TO23 = 0;
parameter signed W38TO24 = 0;
parameter signed W38TO25 = 0;
parameter signed W38TO26 = 0;
parameter signed W38TO27 = 0;
parameter signed W38TO28 = 0;
parameter signed W38TO29 = 0;
parameter signed W38TO30 = 0;
parameter signed W38TO31 = 0;
parameter signed W38TO32 = 0;
parameter signed W38TO33 = 0;
parameter signed W38TO34 = 0;
parameter signed W38TO35 = 0;
parameter signed W38TO36 = 0;
parameter signed W38TO37 = 0;
parameter signed W38TO38 = 0;
parameter signed W38TO39 = 0;
parameter signed W38TO40 = 0;
parameter signed W38TO41 = 0;
parameter signed W38TO42 = 0;
parameter signed W38TO43 = 0;
parameter signed W38TO44 = 0;
parameter signed W38TO45 = 0;
parameter signed W38TO46 = 0;
parameter signed W38TO47 = 0;
parameter signed W38TO48 = 0;
parameter signed W38TO49 = 0;
parameter signed W38TO50 = 0;
parameter signed W38TO51 = 0;
parameter signed W38TO52 = 0;
parameter signed W38TO53 = 0;
parameter signed W38TO54 = 0;
parameter signed W38TO55 = 0;
parameter signed W38TO56 = 0;
parameter signed W38TO57 = 0;
parameter signed W38TO58 = 0;
parameter signed W38TO59 = 0;
parameter signed W38TO60 = 0;
parameter signed W38TO61 = 0;
parameter signed W38TO62 = 0;
parameter signed W38TO63 = 0;
parameter signed W39TO0 = 0;
parameter signed W39TO1 = 0;
parameter signed W39TO2 = 0;
parameter signed W39TO3 = 0;
parameter signed W39TO4 = 0;
parameter signed W39TO5 = 0;
parameter signed W39TO6 = 0;
parameter signed W39TO7 = 0;
parameter signed W39TO8 = 0;
parameter signed W39TO9 = 0;
parameter signed W39TO10 = 0;
parameter signed W39TO11 = 0;
parameter signed W39TO12 = 0;
parameter signed W39TO13 = 0;
parameter signed W39TO14 = 0;
parameter signed W39TO15 = 0;
parameter signed W39TO16 = 0;
parameter signed W39TO17 = 0;
parameter signed W39TO18 = 0;
parameter signed W39TO19 = 0;
parameter signed W39TO20 = 0;
parameter signed W39TO21 = 0;
parameter signed W39TO22 = 0;
parameter signed W39TO23 = 0;
parameter signed W39TO24 = 0;
parameter signed W39TO25 = 0;
parameter signed W39TO26 = 0;
parameter signed W39TO27 = 0;
parameter signed W39TO28 = 0;
parameter signed W39TO29 = 0;
parameter signed W39TO30 = 0;
parameter signed W39TO31 = 0;
parameter signed W39TO32 = 0;
parameter signed W39TO33 = 0;
parameter signed W39TO34 = 0;
parameter signed W39TO35 = 0;
parameter signed W39TO36 = 0;
parameter signed W39TO37 = 0;
parameter signed W39TO38 = 0;
parameter signed W39TO39 = 0;
parameter signed W39TO40 = 0;
parameter signed W39TO41 = 0;
parameter signed W39TO42 = 0;
parameter signed W39TO43 = 0;
parameter signed W39TO44 = 0;
parameter signed W39TO45 = 0;
parameter signed W39TO46 = 0;
parameter signed W39TO47 = 0;
parameter signed W39TO48 = 0;
parameter signed W39TO49 = 0;
parameter signed W39TO50 = 0;
parameter signed W39TO51 = 0;
parameter signed W39TO52 = 0;
parameter signed W39TO53 = 0;
parameter signed W39TO54 = 0;
parameter signed W39TO55 = 0;
parameter signed W39TO56 = 0;
parameter signed W39TO57 = 0;
parameter signed W39TO58 = 0;
parameter signed W39TO59 = 0;
parameter signed W39TO60 = 0;
parameter signed W39TO61 = 0;
parameter signed W39TO62 = 0;
parameter signed W39TO63 = 0;
parameter signed W40TO0 = 0;
parameter signed W40TO1 = 0;
parameter signed W40TO2 = 0;
parameter signed W40TO3 = 0;
parameter signed W40TO4 = 0;
parameter signed W40TO5 = 0;
parameter signed W40TO6 = 0;
parameter signed W40TO7 = 0;
parameter signed W40TO8 = 0;
parameter signed W40TO9 = 0;
parameter signed W40TO10 = 0;
parameter signed W40TO11 = 0;
parameter signed W40TO12 = 0;
parameter signed W40TO13 = 0;
parameter signed W40TO14 = 0;
parameter signed W40TO15 = 0;
parameter signed W40TO16 = 0;
parameter signed W40TO17 = 0;
parameter signed W40TO18 = 0;
parameter signed W40TO19 = 0;
parameter signed W40TO20 = 0;
parameter signed W40TO21 = 0;
parameter signed W40TO22 = 0;
parameter signed W40TO23 = 0;
parameter signed W40TO24 = 0;
parameter signed W40TO25 = 0;
parameter signed W40TO26 = 0;
parameter signed W40TO27 = 0;
parameter signed W40TO28 = 0;
parameter signed W40TO29 = 0;
parameter signed W40TO30 = 0;
parameter signed W40TO31 = 0;
parameter signed W40TO32 = 0;
parameter signed W40TO33 = 0;
parameter signed W40TO34 = 0;
parameter signed W40TO35 = 0;
parameter signed W40TO36 = 0;
parameter signed W40TO37 = 0;
parameter signed W40TO38 = 0;
parameter signed W40TO39 = 0;
parameter signed W40TO40 = 0;
parameter signed W40TO41 = 0;
parameter signed W40TO42 = 0;
parameter signed W40TO43 = 0;
parameter signed W40TO44 = 0;
parameter signed W40TO45 = 0;
parameter signed W40TO46 = 0;
parameter signed W40TO47 = 0;
parameter signed W40TO48 = 0;
parameter signed W40TO49 = 0;
parameter signed W40TO50 = 0;
parameter signed W40TO51 = 0;
parameter signed W40TO52 = 0;
parameter signed W40TO53 = 0;
parameter signed W40TO54 = 0;
parameter signed W40TO55 = 0;
parameter signed W40TO56 = 0;
parameter signed W40TO57 = 0;
parameter signed W40TO58 = 0;
parameter signed W40TO59 = 0;
parameter signed W40TO60 = 0;
parameter signed W40TO61 = 0;
parameter signed W40TO62 = 0;
parameter signed W40TO63 = 0;
parameter signed W41TO0 = 0;
parameter signed W41TO1 = 0;
parameter signed W41TO2 = 0;
parameter signed W41TO3 = 0;
parameter signed W41TO4 = 0;
parameter signed W41TO5 = 0;
parameter signed W41TO6 = 0;
parameter signed W41TO7 = 0;
parameter signed W41TO8 = 0;
parameter signed W41TO9 = 0;
parameter signed W41TO10 = 0;
parameter signed W41TO11 = 0;
parameter signed W41TO12 = 0;
parameter signed W41TO13 = 0;
parameter signed W41TO14 = 0;
parameter signed W41TO15 = 0;
parameter signed W41TO16 = 0;
parameter signed W41TO17 = 0;
parameter signed W41TO18 = 0;
parameter signed W41TO19 = 0;
parameter signed W41TO20 = 0;
parameter signed W41TO21 = 0;
parameter signed W41TO22 = 0;
parameter signed W41TO23 = 0;
parameter signed W41TO24 = 0;
parameter signed W41TO25 = 0;
parameter signed W41TO26 = 0;
parameter signed W41TO27 = 0;
parameter signed W41TO28 = 0;
parameter signed W41TO29 = 0;
parameter signed W41TO30 = 0;
parameter signed W41TO31 = 0;
parameter signed W41TO32 = 0;
parameter signed W41TO33 = 0;
parameter signed W41TO34 = 0;
parameter signed W41TO35 = 0;
parameter signed W41TO36 = 0;
parameter signed W41TO37 = 0;
parameter signed W41TO38 = 0;
parameter signed W41TO39 = 0;
parameter signed W41TO40 = 0;
parameter signed W41TO41 = 0;
parameter signed W41TO42 = 0;
parameter signed W41TO43 = 0;
parameter signed W41TO44 = 0;
parameter signed W41TO45 = 0;
parameter signed W41TO46 = 0;
parameter signed W41TO47 = 0;
parameter signed W41TO48 = 0;
parameter signed W41TO49 = 0;
parameter signed W41TO50 = 0;
parameter signed W41TO51 = 0;
parameter signed W41TO52 = 0;
parameter signed W41TO53 = 0;
parameter signed W41TO54 = 0;
parameter signed W41TO55 = 0;
parameter signed W41TO56 = 0;
parameter signed W41TO57 = 0;
parameter signed W41TO58 = 0;
parameter signed W41TO59 = 0;
parameter signed W41TO60 = 0;
parameter signed W41TO61 = 0;
parameter signed W41TO62 = 0;
parameter signed W41TO63 = 0;
parameter signed W42TO0 = 0;
parameter signed W42TO1 = 0;
parameter signed W42TO2 = 0;
parameter signed W42TO3 = 0;
parameter signed W42TO4 = 0;
parameter signed W42TO5 = 0;
parameter signed W42TO6 = 0;
parameter signed W42TO7 = 0;
parameter signed W42TO8 = 0;
parameter signed W42TO9 = 0;
parameter signed W42TO10 = 0;
parameter signed W42TO11 = 0;
parameter signed W42TO12 = 0;
parameter signed W42TO13 = 0;
parameter signed W42TO14 = 0;
parameter signed W42TO15 = 0;
parameter signed W42TO16 = 0;
parameter signed W42TO17 = 0;
parameter signed W42TO18 = 0;
parameter signed W42TO19 = 0;
parameter signed W42TO20 = 0;
parameter signed W42TO21 = 0;
parameter signed W42TO22 = 0;
parameter signed W42TO23 = 0;
parameter signed W42TO24 = 0;
parameter signed W42TO25 = 0;
parameter signed W42TO26 = 0;
parameter signed W42TO27 = 0;
parameter signed W42TO28 = 0;
parameter signed W42TO29 = 0;
parameter signed W42TO30 = 0;
parameter signed W42TO31 = 0;
parameter signed W42TO32 = 0;
parameter signed W42TO33 = 0;
parameter signed W42TO34 = 0;
parameter signed W42TO35 = 0;
parameter signed W42TO36 = 0;
parameter signed W42TO37 = 0;
parameter signed W42TO38 = 0;
parameter signed W42TO39 = 0;
parameter signed W42TO40 = 0;
parameter signed W42TO41 = 0;
parameter signed W42TO42 = 0;
parameter signed W42TO43 = 0;
parameter signed W42TO44 = 0;
parameter signed W42TO45 = 0;
parameter signed W42TO46 = 0;
parameter signed W42TO47 = 0;
parameter signed W42TO48 = 0;
parameter signed W42TO49 = 0;
parameter signed W42TO50 = 0;
parameter signed W42TO51 = 0;
parameter signed W42TO52 = 0;
parameter signed W42TO53 = 0;
parameter signed W42TO54 = 0;
parameter signed W42TO55 = 0;
parameter signed W42TO56 = 0;
parameter signed W42TO57 = 0;
parameter signed W42TO58 = 0;
parameter signed W42TO59 = 0;
parameter signed W42TO60 = 0;
parameter signed W42TO61 = 0;
parameter signed W42TO62 = 0;
parameter signed W42TO63 = 0;
parameter signed W43TO0 = 0;
parameter signed W43TO1 = 0;
parameter signed W43TO2 = 0;
parameter signed W43TO3 = 0;
parameter signed W43TO4 = 0;
parameter signed W43TO5 = 0;
parameter signed W43TO6 = 0;
parameter signed W43TO7 = 0;
parameter signed W43TO8 = 0;
parameter signed W43TO9 = 0;
parameter signed W43TO10 = 0;
parameter signed W43TO11 = 0;
parameter signed W43TO12 = 0;
parameter signed W43TO13 = 0;
parameter signed W43TO14 = 0;
parameter signed W43TO15 = 0;
parameter signed W43TO16 = 0;
parameter signed W43TO17 = 0;
parameter signed W43TO18 = 0;
parameter signed W43TO19 = 0;
parameter signed W43TO20 = 0;
parameter signed W43TO21 = 0;
parameter signed W43TO22 = 0;
parameter signed W43TO23 = 0;
parameter signed W43TO24 = 0;
parameter signed W43TO25 = 0;
parameter signed W43TO26 = 0;
parameter signed W43TO27 = 0;
parameter signed W43TO28 = 0;
parameter signed W43TO29 = 0;
parameter signed W43TO30 = 0;
parameter signed W43TO31 = 0;
parameter signed W43TO32 = 0;
parameter signed W43TO33 = 0;
parameter signed W43TO34 = 0;
parameter signed W43TO35 = 0;
parameter signed W43TO36 = 0;
parameter signed W43TO37 = 0;
parameter signed W43TO38 = 0;
parameter signed W43TO39 = 0;
parameter signed W43TO40 = 0;
parameter signed W43TO41 = 0;
parameter signed W43TO42 = 0;
parameter signed W43TO43 = 0;
parameter signed W43TO44 = 0;
parameter signed W43TO45 = 0;
parameter signed W43TO46 = 0;
parameter signed W43TO47 = 0;
parameter signed W43TO48 = 0;
parameter signed W43TO49 = 0;
parameter signed W43TO50 = 0;
parameter signed W43TO51 = 0;
parameter signed W43TO52 = 0;
parameter signed W43TO53 = 0;
parameter signed W43TO54 = 0;
parameter signed W43TO55 = 0;
parameter signed W43TO56 = 0;
parameter signed W43TO57 = 0;
parameter signed W43TO58 = 0;
parameter signed W43TO59 = 0;
parameter signed W43TO60 = 0;
parameter signed W43TO61 = 0;
parameter signed W43TO62 = 0;
parameter signed W43TO63 = 0;
parameter signed W44TO0 = 0;
parameter signed W44TO1 = 0;
parameter signed W44TO2 = 0;
parameter signed W44TO3 = 0;
parameter signed W44TO4 = 0;
parameter signed W44TO5 = 0;
parameter signed W44TO6 = 0;
parameter signed W44TO7 = 0;
parameter signed W44TO8 = 0;
parameter signed W44TO9 = 0;
parameter signed W44TO10 = 0;
parameter signed W44TO11 = 0;
parameter signed W44TO12 = 0;
parameter signed W44TO13 = 0;
parameter signed W44TO14 = 0;
parameter signed W44TO15 = 0;
parameter signed W44TO16 = 0;
parameter signed W44TO17 = 0;
parameter signed W44TO18 = 0;
parameter signed W44TO19 = 0;
parameter signed W44TO20 = 0;
parameter signed W44TO21 = 0;
parameter signed W44TO22 = 0;
parameter signed W44TO23 = 0;
parameter signed W44TO24 = 0;
parameter signed W44TO25 = 0;
parameter signed W44TO26 = 0;
parameter signed W44TO27 = 0;
parameter signed W44TO28 = 0;
parameter signed W44TO29 = 0;
parameter signed W44TO30 = 0;
parameter signed W44TO31 = 0;
parameter signed W44TO32 = 0;
parameter signed W44TO33 = 0;
parameter signed W44TO34 = 0;
parameter signed W44TO35 = 0;
parameter signed W44TO36 = 0;
parameter signed W44TO37 = 0;
parameter signed W44TO38 = 0;
parameter signed W44TO39 = 0;
parameter signed W44TO40 = 0;
parameter signed W44TO41 = 0;
parameter signed W44TO42 = 0;
parameter signed W44TO43 = 0;
parameter signed W44TO44 = 0;
parameter signed W44TO45 = 0;
parameter signed W44TO46 = 0;
parameter signed W44TO47 = 0;
parameter signed W44TO48 = 0;
parameter signed W44TO49 = 0;
parameter signed W44TO50 = 0;
parameter signed W44TO51 = 0;
parameter signed W44TO52 = 0;
parameter signed W44TO53 = 0;
parameter signed W44TO54 = 0;
parameter signed W44TO55 = 0;
parameter signed W44TO56 = 0;
parameter signed W44TO57 = 0;
parameter signed W44TO58 = 0;
parameter signed W44TO59 = 0;
parameter signed W44TO60 = 0;
parameter signed W44TO61 = 0;
parameter signed W44TO62 = 0;
parameter signed W44TO63 = 0;
parameter signed W45TO0 = 0;
parameter signed W45TO1 = 0;
parameter signed W45TO2 = 0;
parameter signed W45TO3 = 0;
parameter signed W45TO4 = 0;
parameter signed W45TO5 = 0;
parameter signed W45TO6 = 0;
parameter signed W45TO7 = 0;
parameter signed W45TO8 = 0;
parameter signed W45TO9 = 0;
parameter signed W45TO10 = 0;
parameter signed W45TO11 = 0;
parameter signed W45TO12 = 0;
parameter signed W45TO13 = 0;
parameter signed W45TO14 = 0;
parameter signed W45TO15 = 0;
parameter signed W45TO16 = 0;
parameter signed W45TO17 = 0;
parameter signed W45TO18 = 0;
parameter signed W45TO19 = 0;
parameter signed W45TO20 = 0;
parameter signed W45TO21 = 0;
parameter signed W45TO22 = 0;
parameter signed W45TO23 = 0;
parameter signed W45TO24 = 0;
parameter signed W45TO25 = 0;
parameter signed W45TO26 = 0;
parameter signed W45TO27 = 0;
parameter signed W45TO28 = 0;
parameter signed W45TO29 = 0;
parameter signed W45TO30 = 0;
parameter signed W45TO31 = 0;
parameter signed W45TO32 = 0;
parameter signed W45TO33 = 0;
parameter signed W45TO34 = 0;
parameter signed W45TO35 = 0;
parameter signed W45TO36 = 0;
parameter signed W45TO37 = 0;
parameter signed W45TO38 = 0;
parameter signed W45TO39 = 0;
parameter signed W45TO40 = 0;
parameter signed W45TO41 = 0;
parameter signed W45TO42 = 0;
parameter signed W45TO43 = 0;
parameter signed W45TO44 = 0;
parameter signed W45TO45 = 0;
parameter signed W45TO46 = 0;
parameter signed W45TO47 = 0;
parameter signed W45TO48 = 0;
parameter signed W45TO49 = 0;
parameter signed W45TO50 = 0;
parameter signed W45TO51 = 0;
parameter signed W45TO52 = 0;
parameter signed W45TO53 = 0;
parameter signed W45TO54 = 0;
parameter signed W45TO55 = 0;
parameter signed W45TO56 = 0;
parameter signed W45TO57 = 0;
parameter signed W45TO58 = 0;
parameter signed W45TO59 = 0;
parameter signed W45TO60 = 0;
parameter signed W45TO61 = 0;
parameter signed W45TO62 = 0;
parameter signed W45TO63 = 0;
parameter signed W46TO0 = 0;
parameter signed W46TO1 = 0;
parameter signed W46TO2 = 0;
parameter signed W46TO3 = 0;
parameter signed W46TO4 = 0;
parameter signed W46TO5 = 0;
parameter signed W46TO6 = 0;
parameter signed W46TO7 = 0;
parameter signed W46TO8 = 0;
parameter signed W46TO9 = 0;
parameter signed W46TO10 = 0;
parameter signed W46TO11 = 0;
parameter signed W46TO12 = 0;
parameter signed W46TO13 = 0;
parameter signed W46TO14 = 0;
parameter signed W46TO15 = 0;
parameter signed W46TO16 = 0;
parameter signed W46TO17 = 0;
parameter signed W46TO18 = 0;
parameter signed W46TO19 = 0;
parameter signed W46TO20 = 0;
parameter signed W46TO21 = 0;
parameter signed W46TO22 = 0;
parameter signed W46TO23 = 0;
parameter signed W46TO24 = 0;
parameter signed W46TO25 = 0;
parameter signed W46TO26 = 0;
parameter signed W46TO27 = 0;
parameter signed W46TO28 = 0;
parameter signed W46TO29 = 0;
parameter signed W46TO30 = 0;
parameter signed W46TO31 = 0;
parameter signed W46TO32 = 0;
parameter signed W46TO33 = 0;
parameter signed W46TO34 = 0;
parameter signed W46TO35 = 0;
parameter signed W46TO36 = 0;
parameter signed W46TO37 = 0;
parameter signed W46TO38 = 0;
parameter signed W46TO39 = 0;
parameter signed W46TO40 = 0;
parameter signed W46TO41 = 0;
parameter signed W46TO42 = 0;
parameter signed W46TO43 = 0;
parameter signed W46TO44 = 0;
parameter signed W46TO45 = 0;
parameter signed W46TO46 = 0;
parameter signed W46TO47 = 0;
parameter signed W46TO48 = 0;
parameter signed W46TO49 = 0;
parameter signed W46TO50 = 0;
parameter signed W46TO51 = 0;
parameter signed W46TO52 = 0;
parameter signed W46TO53 = 0;
parameter signed W46TO54 = 0;
parameter signed W46TO55 = 0;
parameter signed W46TO56 = 0;
parameter signed W46TO57 = 0;
parameter signed W46TO58 = 0;
parameter signed W46TO59 = 0;
parameter signed W46TO60 = 0;
parameter signed W46TO61 = 0;
parameter signed W46TO62 = 0;
parameter signed W46TO63 = 0;
parameter signed W47TO0 = 0;
parameter signed W47TO1 = 0;
parameter signed W47TO2 = 0;
parameter signed W47TO3 = 0;
parameter signed W47TO4 = 0;
parameter signed W47TO5 = 0;
parameter signed W47TO6 = 0;
parameter signed W47TO7 = 0;
parameter signed W47TO8 = 0;
parameter signed W47TO9 = 0;
parameter signed W47TO10 = 0;
parameter signed W47TO11 = 0;
parameter signed W47TO12 = 0;
parameter signed W47TO13 = 0;
parameter signed W47TO14 = 0;
parameter signed W47TO15 = 0;
parameter signed W47TO16 = 0;
parameter signed W47TO17 = 0;
parameter signed W47TO18 = 0;
parameter signed W47TO19 = 0;
parameter signed W47TO20 = 0;
parameter signed W47TO21 = 0;
parameter signed W47TO22 = 0;
parameter signed W47TO23 = 0;
parameter signed W47TO24 = 0;
parameter signed W47TO25 = 0;
parameter signed W47TO26 = 0;
parameter signed W47TO27 = 0;
parameter signed W47TO28 = 0;
parameter signed W47TO29 = 0;
parameter signed W47TO30 = 0;
parameter signed W47TO31 = 0;
parameter signed W47TO32 = 0;
parameter signed W47TO33 = 0;
parameter signed W47TO34 = 0;
parameter signed W47TO35 = 0;
parameter signed W47TO36 = 0;
parameter signed W47TO37 = 0;
parameter signed W47TO38 = 0;
parameter signed W47TO39 = 0;
parameter signed W47TO40 = 0;
parameter signed W47TO41 = 0;
parameter signed W47TO42 = 0;
parameter signed W47TO43 = 0;
parameter signed W47TO44 = 0;
parameter signed W47TO45 = 0;
parameter signed W47TO46 = 0;
parameter signed W47TO47 = 0;
parameter signed W47TO48 = 0;
parameter signed W47TO49 = 0;
parameter signed W47TO50 = 0;
parameter signed W47TO51 = 0;
parameter signed W47TO52 = 0;
parameter signed W47TO53 = 0;
parameter signed W47TO54 = 0;
parameter signed W47TO55 = 0;
parameter signed W47TO56 = 0;
parameter signed W47TO57 = 0;
parameter signed W47TO58 = 0;
parameter signed W47TO59 = 0;
parameter signed W47TO60 = 0;
parameter signed W47TO61 = 0;
parameter signed W47TO62 = 0;
parameter signed W47TO63 = 0;
parameter signed W48TO0 = 0;
parameter signed W48TO1 = 0;
parameter signed W48TO2 = 0;
parameter signed W48TO3 = 0;
parameter signed W48TO4 = 0;
parameter signed W48TO5 = 0;
parameter signed W48TO6 = 0;
parameter signed W48TO7 = 0;
parameter signed W48TO8 = 0;
parameter signed W48TO9 = 0;
parameter signed W48TO10 = 0;
parameter signed W48TO11 = 0;
parameter signed W48TO12 = 0;
parameter signed W48TO13 = 0;
parameter signed W48TO14 = 0;
parameter signed W48TO15 = 0;
parameter signed W48TO16 = 0;
parameter signed W48TO17 = 0;
parameter signed W48TO18 = 0;
parameter signed W48TO19 = 0;
parameter signed W48TO20 = 0;
parameter signed W48TO21 = 0;
parameter signed W48TO22 = 0;
parameter signed W48TO23 = 0;
parameter signed W48TO24 = 0;
parameter signed W48TO25 = 0;
parameter signed W48TO26 = 0;
parameter signed W48TO27 = 0;
parameter signed W48TO28 = 0;
parameter signed W48TO29 = 0;
parameter signed W48TO30 = 0;
parameter signed W48TO31 = 0;
parameter signed W48TO32 = 0;
parameter signed W48TO33 = 0;
parameter signed W48TO34 = 0;
parameter signed W48TO35 = 0;
parameter signed W48TO36 = 0;
parameter signed W48TO37 = 0;
parameter signed W48TO38 = 0;
parameter signed W48TO39 = 0;
parameter signed W48TO40 = 0;
parameter signed W48TO41 = 0;
parameter signed W48TO42 = 0;
parameter signed W48TO43 = 0;
parameter signed W48TO44 = 0;
parameter signed W48TO45 = 0;
parameter signed W48TO46 = 0;
parameter signed W48TO47 = 0;
parameter signed W48TO48 = 0;
parameter signed W48TO49 = 0;
parameter signed W48TO50 = 0;
parameter signed W48TO51 = 0;
parameter signed W48TO52 = 0;
parameter signed W48TO53 = 0;
parameter signed W48TO54 = 0;
parameter signed W48TO55 = 0;
parameter signed W48TO56 = 0;
parameter signed W48TO57 = 0;
parameter signed W48TO58 = 0;
parameter signed W48TO59 = 0;
parameter signed W48TO60 = 0;
parameter signed W48TO61 = 0;
parameter signed W48TO62 = 0;
parameter signed W48TO63 = 0;
parameter signed W49TO0 = 0;
parameter signed W49TO1 = 0;
parameter signed W49TO2 = 0;
parameter signed W49TO3 = 0;
parameter signed W49TO4 = 0;
parameter signed W49TO5 = 0;
parameter signed W49TO6 = 0;
parameter signed W49TO7 = 0;
parameter signed W49TO8 = 0;
parameter signed W49TO9 = 0;
parameter signed W49TO10 = 0;
parameter signed W49TO11 = 0;
parameter signed W49TO12 = 0;
parameter signed W49TO13 = 0;
parameter signed W49TO14 = 0;
parameter signed W49TO15 = 0;
parameter signed W49TO16 = 0;
parameter signed W49TO17 = 0;
parameter signed W49TO18 = 0;
parameter signed W49TO19 = 0;
parameter signed W49TO20 = 0;
parameter signed W49TO21 = 0;
parameter signed W49TO22 = 0;
parameter signed W49TO23 = 0;
parameter signed W49TO24 = 0;
parameter signed W49TO25 = 0;
parameter signed W49TO26 = 0;
parameter signed W49TO27 = 0;
parameter signed W49TO28 = 0;
parameter signed W49TO29 = 0;
parameter signed W49TO30 = 0;
parameter signed W49TO31 = 0;
parameter signed W49TO32 = 0;
parameter signed W49TO33 = 0;
parameter signed W49TO34 = 0;
parameter signed W49TO35 = 0;
parameter signed W49TO36 = 0;
parameter signed W49TO37 = 0;
parameter signed W49TO38 = 0;
parameter signed W49TO39 = 0;
parameter signed W49TO40 = 0;
parameter signed W49TO41 = 0;
parameter signed W49TO42 = 0;
parameter signed W49TO43 = 0;
parameter signed W49TO44 = 0;
parameter signed W49TO45 = 0;
parameter signed W49TO46 = 0;
parameter signed W49TO47 = 0;
parameter signed W49TO48 = 0;
parameter signed W49TO49 = 0;
parameter signed W49TO50 = 0;
parameter signed W49TO51 = 0;
parameter signed W49TO52 = 0;
parameter signed W49TO53 = 0;
parameter signed W49TO54 = 0;
parameter signed W49TO55 = 0;
parameter signed W49TO56 = 0;
parameter signed W49TO57 = 0;
parameter signed W49TO58 = 0;
parameter signed W49TO59 = 0;
parameter signed W49TO60 = 0;
parameter signed W49TO61 = 0;
parameter signed W49TO62 = 0;
parameter signed W49TO63 = 0;
parameter signed W50TO0 = 0;
parameter signed W50TO1 = 0;
parameter signed W50TO2 = 0;
parameter signed W50TO3 = 0;
parameter signed W50TO4 = 0;
parameter signed W50TO5 = 0;
parameter signed W50TO6 = 0;
parameter signed W50TO7 = 0;
parameter signed W50TO8 = 0;
parameter signed W50TO9 = 0;
parameter signed W50TO10 = 0;
parameter signed W50TO11 = 0;
parameter signed W50TO12 = 0;
parameter signed W50TO13 = 0;
parameter signed W50TO14 = 0;
parameter signed W50TO15 = 0;
parameter signed W50TO16 = 0;
parameter signed W50TO17 = 0;
parameter signed W50TO18 = 0;
parameter signed W50TO19 = 0;
parameter signed W50TO20 = 0;
parameter signed W50TO21 = 0;
parameter signed W50TO22 = 0;
parameter signed W50TO23 = 0;
parameter signed W50TO24 = 0;
parameter signed W50TO25 = 0;
parameter signed W50TO26 = 0;
parameter signed W50TO27 = 0;
parameter signed W50TO28 = 0;
parameter signed W50TO29 = 0;
parameter signed W50TO30 = 0;
parameter signed W50TO31 = 0;
parameter signed W50TO32 = 0;
parameter signed W50TO33 = 0;
parameter signed W50TO34 = 0;
parameter signed W50TO35 = 0;
parameter signed W50TO36 = 0;
parameter signed W50TO37 = 0;
parameter signed W50TO38 = 0;
parameter signed W50TO39 = 0;
parameter signed W50TO40 = 0;
parameter signed W50TO41 = 0;
parameter signed W50TO42 = 0;
parameter signed W50TO43 = 0;
parameter signed W50TO44 = 0;
parameter signed W50TO45 = 0;
parameter signed W50TO46 = 0;
parameter signed W50TO47 = 0;
parameter signed W50TO48 = 0;
parameter signed W50TO49 = 0;
parameter signed W50TO50 = 0;
parameter signed W50TO51 = 0;
parameter signed W50TO52 = 0;
parameter signed W50TO53 = 0;
parameter signed W50TO54 = 0;
parameter signed W50TO55 = 0;
parameter signed W50TO56 = 0;
parameter signed W50TO57 = 0;
parameter signed W50TO58 = 0;
parameter signed W50TO59 = 0;
parameter signed W50TO60 = 0;
parameter signed W50TO61 = 0;
parameter signed W50TO62 = 0;
parameter signed W50TO63 = 0;
parameter signed W51TO0 = 0;
parameter signed W51TO1 = 0;
parameter signed W51TO2 = 0;
parameter signed W51TO3 = 0;
parameter signed W51TO4 = 0;
parameter signed W51TO5 = 0;
parameter signed W51TO6 = 0;
parameter signed W51TO7 = 0;
parameter signed W51TO8 = 0;
parameter signed W51TO9 = 0;
parameter signed W51TO10 = 0;
parameter signed W51TO11 = 0;
parameter signed W51TO12 = 0;
parameter signed W51TO13 = 0;
parameter signed W51TO14 = 0;
parameter signed W51TO15 = 0;
parameter signed W51TO16 = 0;
parameter signed W51TO17 = 0;
parameter signed W51TO18 = 0;
parameter signed W51TO19 = 0;
parameter signed W51TO20 = 0;
parameter signed W51TO21 = 0;
parameter signed W51TO22 = 0;
parameter signed W51TO23 = 0;
parameter signed W51TO24 = 0;
parameter signed W51TO25 = 0;
parameter signed W51TO26 = 0;
parameter signed W51TO27 = 0;
parameter signed W51TO28 = 0;
parameter signed W51TO29 = 0;
parameter signed W51TO30 = 0;
parameter signed W51TO31 = 0;
parameter signed W51TO32 = 0;
parameter signed W51TO33 = 0;
parameter signed W51TO34 = 0;
parameter signed W51TO35 = 0;
parameter signed W51TO36 = 0;
parameter signed W51TO37 = 0;
parameter signed W51TO38 = 0;
parameter signed W51TO39 = 0;
parameter signed W51TO40 = 0;
parameter signed W51TO41 = 0;
parameter signed W51TO42 = 0;
parameter signed W51TO43 = 0;
parameter signed W51TO44 = 0;
parameter signed W51TO45 = 0;
parameter signed W51TO46 = 0;
parameter signed W51TO47 = 0;
parameter signed W51TO48 = 0;
parameter signed W51TO49 = 0;
parameter signed W51TO50 = 0;
parameter signed W51TO51 = 0;
parameter signed W51TO52 = 0;
parameter signed W51TO53 = 0;
parameter signed W51TO54 = 0;
parameter signed W51TO55 = 0;
parameter signed W51TO56 = 0;
parameter signed W51TO57 = 0;
parameter signed W51TO58 = 0;
parameter signed W51TO59 = 0;
parameter signed W51TO60 = 0;
parameter signed W51TO61 = 0;
parameter signed W51TO62 = 0;
parameter signed W51TO63 = 0;
parameter signed W52TO0 = 0;
parameter signed W52TO1 = 0;
parameter signed W52TO2 = 0;
parameter signed W52TO3 = 0;
parameter signed W52TO4 = 0;
parameter signed W52TO5 = 0;
parameter signed W52TO6 = 0;
parameter signed W52TO7 = 0;
parameter signed W52TO8 = 0;
parameter signed W52TO9 = 0;
parameter signed W52TO10 = 0;
parameter signed W52TO11 = 0;
parameter signed W52TO12 = 0;
parameter signed W52TO13 = 0;
parameter signed W52TO14 = 0;
parameter signed W52TO15 = 0;
parameter signed W52TO16 = 0;
parameter signed W52TO17 = 0;
parameter signed W52TO18 = 0;
parameter signed W52TO19 = 0;
parameter signed W52TO20 = 0;
parameter signed W52TO21 = 0;
parameter signed W52TO22 = 0;
parameter signed W52TO23 = 0;
parameter signed W52TO24 = 0;
parameter signed W52TO25 = 0;
parameter signed W52TO26 = 0;
parameter signed W52TO27 = 0;
parameter signed W52TO28 = 0;
parameter signed W52TO29 = 0;
parameter signed W52TO30 = 0;
parameter signed W52TO31 = 0;
parameter signed W52TO32 = 0;
parameter signed W52TO33 = 0;
parameter signed W52TO34 = 0;
parameter signed W52TO35 = 0;
parameter signed W52TO36 = 0;
parameter signed W52TO37 = 0;
parameter signed W52TO38 = 0;
parameter signed W52TO39 = 0;
parameter signed W52TO40 = 0;
parameter signed W52TO41 = 0;
parameter signed W52TO42 = 0;
parameter signed W52TO43 = 0;
parameter signed W52TO44 = 0;
parameter signed W52TO45 = 0;
parameter signed W52TO46 = 0;
parameter signed W52TO47 = 0;
parameter signed W52TO48 = 0;
parameter signed W52TO49 = 0;
parameter signed W52TO50 = 0;
parameter signed W52TO51 = 0;
parameter signed W52TO52 = 0;
parameter signed W52TO53 = 0;
parameter signed W52TO54 = 0;
parameter signed W52TO55 = 0;
parameter signed W52TO56 = 0;
parameter signed W52TO57 = 0;
parameter signed W52TO58 = 0;
parameter signed W52TO59 = 0;
parameter signed W52TO60 = 0;
parameter signed W52TO61 = 0;
parameter signed W52TO62 = 0;
parameter signed W52TO63 = 0;
parameter signed W53TO0 = 0;
parameter signed W53TO1 = 0;
parameter signed W53TO2 = 0;
parameter signed W53TO3 = 0;
parameter signed W53TO4 = 0;
parameter signed W53TO5 = 0;
parameter signed W53TO6 = 0;
parameter signed W53TO7 = 0;
parameter signed W53TO8 = 0;
parameter signed W53TO9 = 0;
parameter signed W53TO10 = 0;
parameter signed W53TO11 = 0;
parameter signed W53TO12 = 0;
parameter signed W53TO13 = 0;
parameter signed W53TO14 = 0;
parameter signed W53TO15 = 0;
parameter signed W53TO16 = 0;
parameter signed W53TO17 = 0;
parameter signed W53TO18 = 0;
parameter signed W53TO19 = 0;
parameter signed W53TO20 = 0;
parameter signed W53TO21 = 0;
parameter signed W53TO22 = 0;
parameter signed W53TO23 = 0;
parameter signed W53TO24 = 0;
parameter signed W53TO25 = 0;
parameter signed W53TO26 = 0;
parameter signed W53TO27 = 0;
parameter signed W53TO28 = 0;
parameter signed W53TO29 = 0;
parameter signed W53TO30 = 0;
parameter signed W53TO31 = 0;
parameter signed W53TO32 = 0;
parameter signed W53TO33 = 0;
parameter signed W53TO34 = 0;
parameter signed W53TO35 = 0;
parameter signed W53TO36 = 0;
parameter signed W53TO37 = 0;
parameter signed W53TO38 = 0;
parameter signed W53TO39 = 0;
parameter signed W53TO40 = 0;
parameter signed W53TO41 = 0;
parameter signed W53TO42 = 0;
parameter signed W53TO43 = 0;
parameter signed W53TO44 = 0;
parameter signed W53TO45 = 0;
parameter signed W53TO46 = 0;
parameter signed W53TO47 = 0;
parameter signed W53TO48 = 0;
parameter signed W53TO49 = 0;
parameter signed W53TO50 = 0;
parameter signed W53TO51 = 0;
parameter signed W53TO52 = 0;
parameter signed W53TO53 = 0;
parameter signed W53TO54 = 0;
parameter signed W53TO55 = 0;
parameter signed W53TO56 = 0;
parameter signed W53TO57 = 0;
parameter signed W53TO58 = 0;
parameter signed W53TO59 = 0;
parameter signed W53TO60 = 0;
parameter signed W53TO61 = 0;
parameter signed W53TO62 = 0;
parameter signed W53TO63 = 0;
parameter signed W54TO0 = 0;
parameter signed W54TO1 = 0;
parameter signed W54TO2 = 0;
parameter signed W54TO3 = 0;
parameter signed W54TO4 = 0;
parameter signed W54TO5 = 0;
parameter signed W54TO6 = 0;
parameter signed W54TO7 = 0;
parameter signed W54TO8 = 0;
parameter signed W54TO9 = 0;
parameter signed W54TO10 = 0;
parameter signed W54TO11 = 0;
parameter signed W54TO12 = 0;
parameter signed W54TO13 = 0;
parameter signed W54TO14 = 0;
parameter signed W54TO15 = 0;
parameter signed W54TO16 = 0;
parameter signed W54TO17 = 0;
parameter signed W54TO18 = 0;
parameter signed W54TO19 = 0;
parameter signed W54TO20 = 0;
parameter signed W54TO21 = 0;
parameter signed W54TO22 = 0;
parameter signed W54TO23 = 0;
parameter signed W54TO24 = 0;
parameter signed W54TO25 = 0;
parameter signed W54TO26 = 0;
parameter signed W54TO27 = 0;
parameter signed W54TO28 = 0;
parameter signed W54TO29 = 0;
parameter signed W54TO30 = 0;
parameter signed W54TO31 = 0;
parameter signed W54TO32 = 0;
parameter signed W54TO33 = 0;
parameter signed W54TO34 = 0;
parameter signed W54TO35 = 0;
parameter signed W54TO36 = 0;
parameter signed W54TO37 = 0;
parameter signed W54TO38 = 0;
parameter signed W54TO39 = 0;
parameter signed W54TO40 = 0;
parameter signed W54TO41 = 0;
parameter signed W54TO42 = 0;
parameter signed W54TO43 = 0;
parameter signed W54TO44 = 0;
parameter signed W54TO45 = 0;
parameter signed W54TO46 = 0;
parameter signed W54TO47 = 0;
parameter signed W54TO48 = 0;
parameter signed W54TO49 = 0;
parameter signed W54TO50 = 0;
parameter signed W54TO51 = 0;
parameter signed W54TO52 = 0;
parameter signed W54TO53 = 0;
parameter signed W54TO54 = 0;
parameter signed W54TO55 = 0;
parameter signed W54TO56 = 0;
parameter signed W54TO57 = 0;
parameter signed W54TO58 = 0;
parameter signed W54TO59 = 0;
parameter signed W54TO60 = 0;
parameter signed W54TO61 = 0;
parameter signed W54TO62 = 0;
parameter signed W54TO63 = 0;
parameter signed W55TO0 = 0;
parameter signed W55TO1 = 0;
parameter signed W55TO2 = 0;
parameter signed W55TO3 = 0;
parameter signed W55TO4 = 0;
parameter signed W55TO5 = 0;
parameter signed W55TO6 = 0;
parameter signed W55TO7 = 0;
parameter signed W55TO8 = 0;
parameter signed W55TO9 = 0;
parameter signed W55TO10 = 0;
parameter signed W55TO11 = 0;
parameter signed W55TO12 = 0;
parameter signed W55TO13 = 0;
parameter signed W55TO14 = 0;
parameter signed W55TO15 = 0;
parameter signed W55TO16 = 0;
parameter signed W55TO17 = 0;
parameter signed W55TO18 = 0;
parameter signed W55TO19 = 0;
parameter signed W55TO20 = 0;
parameter signed W55TO21 = 0;
parameter signed W55TO22 = 0;
parameter signed W55TO23 = 0;
parameter signed W55TO24 = 0;
parameter signed W55TO25 = 0;
parameter signed W55TO26 = 0;
parameter signed W55TO27 = 0;
parameter signed W55TO28 = 0;
parameter signed W55TO29 = 0;
parameter signed W55TO30 = 0;
parameter signed W55TO31 = 0;
parameter signed W55TO32 = 0;
parameter signed W55TO33 = 0;
parameter signed W55TO34 = 0;
parameter signed W55TO35 = 0;
parameter signed W55TO36 = 0;
parameter signed W55TO37 = 0;
parameter signed W55TO38 = 0;
parameter signed W55TO39 = 0;
parameter signed W55TO40 = 0;
parameter signed W55TO41 = 0;
parameter signed W55TO42 = 0;
parameter signed W55TO43 = 0;
parameter signed W55TO44 = 0;
parameter signed W55TO45 = 0;
parameter signed W55TO46 = 0;
parameter signed W55TO47 = 0;
parameter signed W55TO48 = 0;
parameter signed W55TO49 = 0;
parameter signed W55TO50 = 0;
parameter signed W55TO51 = 0;
parameter signed W55TO52 = 0;
parameter signed W55TO53 = 0;
parameter signed W55TO54 = 0;
parameter signed W55TO55 = 0;
parameter signed W55TO56 = 0;
parameter signed W55TO57 = 0;
parameter signed W55TO58 = 0;
parameter signed W55TO59 = 0;
parameter signed W55TO60 = 0;
parameter signed W55TO61 = 0;
parameter signed W55TO62 = 0;
parameter signed W55TO63 = 0;
parameter signed W56TO0 = 0;
parameter signed W56TO1 = 0;
parameter signed W56TO2 = 0;
parameter signed W56TO3 = 0;
parameter signed W56TO4 = 0;
parameter signed W56TO5 = 0;
parameter signed W56TO6 = 0;
parameter signed W56TO7 = 0;
parameter signed W56TO8 = 0;
parameter signed W56TO9 = 0;
parameter signed W56TO10 = 0;
parameter signed W56TO11 = 0;
parameter signed W56TO12 = 0;
parameter signed W56TO13 = 0;
parameter signed W56TO14 = 0;
parameter signed W56TO15 = 0;
parameter signed W56TO16 = 0;
parameter signed W56TO17 = 0;
parameter signed W56TO18 = 0;
parameter signed W56TO19 = 0;
parameter signed W56TO20 = 0;
parameter signed W56TO21 = 0;
parameter signed W56TO22 = 0;
parameter signed W56TO23 = 0;
parameter signed W56TO24 = 0;
parameter signed W56TO25 = 0;
parameter signed W56TO26 = 0;
parameter signed W56TO27 = 0;
parameter signed W56TO28 = 0;
parameter signed W56TO29 = 0;
parameter signed W56TO30 = 0;
parameter signed W56TO31 = 0;
parameter signed W56TO32 = 0;
parameter signed W56TO33 = 0;
parameter signed W56TO34 = 0;
parameter signed W56TO35 = 0;
parameter signed W56TO36 = 0;
parameter signed W56TO37 = 0;
parameter signed W56TO38 = 0;
parameter signed W56TO39 = 0;
parameter signed W56TO40 = 0;
parameter signed W56TO41 = 0;
parameter signed W56TO42 = 0;
parameter signed W56TO43 = 0;
parameter signed W56TO44 = 0;
parameter signed W56TO45 = 0;
parameter signed W56TO46 = 0;
parameter signed W56TO47 = 0;
parameter signed W56TO48 = 0;
parameter signed W56TO49 = 0;
parameter signed W56TO50 = 0;
parameter signed W56TO51 = 0;
parameter signed W56TO52 = 0;
parameter signed W56TO53 = 0;
parameter signed W56TO54 = 0;
parameter signed W56TO55 = 0;
parameter signed W56TO56 = 0;
parameter signed W56TO57 = 0;
parameter signed W56TO58 = 0;
parameter signed W56TO59 = 0;
parameter signed W56TO60 = 0;
parameter signed W56TO61 = 0;
parameter signed W56TO62 = 0;
parameter signed W56TO63 = 0;
parameter signed W57TO0 = 0;
parameter signed W57TO1 = 0;
parameter signed W57TO2 = 0;
parameter signed W57TO3 = 0;
parameter signed W57TO4 = 0;
parameter signed W57TO5 = 0;
parameter signed W57TO6 = 0;
parameter signed W57TO7 = 0;
parameter signed W57TO8 = 0;
parameter signed W57TO9 = 0;
parameter signed W57TO10 = 0;
parameter signed W57TO11 = 0;
parameter signed W57TO12 = 0;
parameter signed W57TO13 = 0;
parameter signed W57TO14 = 0;
parameter signed W57TO15 = 0;
parameter signed W57TO16 = 0;
parameter signed W57TO17 = 0;
parameter signed W57TO18 = 0;
parameter signed W57TO19 = 0;
parameter signed W57TO20 = 0;
parameter signed W57TO21 = 0;
parameter signed W57TO22 = 0;
parameter signed W57TO23 = 0;
parameter signed W57TO24 = 0;
parameter signed W57TO25 = 0;
parameter signed W57TO26 = 0;
parameter signed W57TO27 = 0;
parameter signed W57TO28 = 0;
parameter signed W57TO29 = 0;
parameter signed W57TO30 = 0;
parameter signed W57TO31 = 0;
parameter signed W57TO32 = 0;
parameter signed W57TO33 = 0;
parameter signed W57TO34 = 0;
parameter signed W57TO35 = 0;
parameter signed W57TO36 = 0;
parameter signed W57TO37 = 0;
parameter signed W57TO38 = 0;
parameter signed W57TO39 = 0;
parameter signed W57TO40 = 0;
parameter signed W57TO41 = 0;
parameter signed W57TO42 = 0;
parameter signed W57TO43 = 0;
parameter signed W57TO44 = 0;
parameter signed W57TO45 = 0;
parameter signed W57TO46 = 0;
parameter signed W57TO47 = 0;
parameter signed W57TO48 = 0;
parameter signed W57TO49 = 0;
parameter signed W57TO50 = 0;
parameter signed W57TO51 = 0;
parameter signed W57TO52 = 0;
parameter signed W57TO53 = 0;
parameter signed W57TO54 = 0;
parameter signed W57TO55 = 0;
parameter signed W57TO56 = 0;
parameter signed W57TO57 = 0;
parameter signed W57TO58 = 0;
parameter signed W57TO59 = 0;
parameter signed W57TO60 = 0;
parameter signed W57TO61 = 0;
parameter signed W57TO62 = 0;
parameter signed W57TO63 = 0;
parameter signed W58TO0 = 0;
parameter signed W58TO1 = 0;
parameter signed W58TO2 = 0;
parameter signed W58TO3 = 0;
parameter signed W58TO4 = 0;
parameter signed W58TO5 = 0;
parameter signed W58TO6 = 0;
parameter signed W58TO7 = 0;
parameter signed W58TO8 = 0;
parameter signed W58TO9 = 0;
parameter signed W58TO10 = 0;
parameter signed W58TO11 = 0;
parameter signed W58TO12 = 0;
parameter signed W58TO13 = 0;
parameter signed W58TO14 = 0;
parameter signed W58TO15 = 0;
parameter signed W58TO16 = 0;
parameter signed W58TO17 = 0;
parameter signed W58TO18 = 0;
parameter signed W58TO19 = 0;
parameter signed W58TO20 = 0;
parameter signed W58TO21 = 0;
parameter signed W58TO22 = 0;
parameter signed W58TO23 = 0;
parameter signed W58TO24 = 0;
parameter signed W58TO25 = 0;
parameter signed W58TO26 = 0;
parameter signed W58TO27 = 0;
parameter signed W58TO28 = 0;
parameter signed W58TO29 = 0;
parameter signed W58TO30 = 0;
parameter signed W58TO31 = 0;
parameter signed W58TO32 = 0;
parameter signed W58TO33 = 0;
parameter signed W58TO34 = 0;
parameter signed W58TO35 = 0;
parameter signed W58TO36 = 0;
parameter signed W58TO37 = 0;
parameter signed W58TO38 = 0;
parameter signed W58TO39 = 0;
parameter signed W58TO40 = 0;
parameter signed W58TO41 = 0;
parameter signed W58TO42 = 0;
parameter signed W58TO43 = 0;
parameter signed W58TO44 = 0;
parameter signed W58TO45 = 0;
parameter signed W58TO46 = 0;
parameter signed W58TO47 = 0;
parameter signed W58TO48 = 0;
parameter signed W58TO49 = 0;
parameter signed W58TO50 = 0;
parameter signed W58TO51 = 0;
parameter signed W58TO52 = 0;
parameter signed W58TO53 = 0;
parameter signed W58TO54 = 0;
parameter signed W58TO55 = 0;
parameter signed W58TO56 = 0;
parameter signed W58TO57 = 0;
parameter signed W58TO58 = 0;
parameter signed W58TO59 = 0;
parameter signed W58TO60 = 0;
parameter signed W58TO61 = 0;
parameter signed W58TO62 = 0;
parameter signed W58TO63 = 0;
parameter signed W59TO0 = 0;
parameter signed W59TO1 = 0;
parameter signed W59TO2 = 0;
parameter signed W59TO3 = 0;
parameter signed W59TO4 = 0;
parameter signed W59TO5 = 0;
parameter signed W59TO6 = 0;
parameter signed W59TO7 = 0;
parameter signed W59TO8 = 0;
parameter signed W59TO9 = 0;
parameter signed W59TO10 = 0;
parameter signed W59TO11 = 0;
parameter signed W59TO12 = 0;
parameter signed W59TO13 = 0;
parameter signed W59TO14 = 0;
parameter signed W59TO15 = 0;
parameter signed W59TO16 = 0;
parameter signed W59TO17 = 0;
parameter signed W59TO18 = 0;
parameter signed W59TO19 = 0;
parameter signed W59TO20 = 0;
parameter signed W59TO21 = 0;
parameter signed W59TO22 = 0;
parameter signed W59TO23 = 0;
parameter signed W59TO24 = 0;
parameter signed W59TO25 = 0;
parameter signed W59TO26 = 0;
parameter signed W59TO27 = 0;
parameter signed W59TO28 = 0;
parameter signed W59TO29 = 0;
parameter signed W59TO30 = 0;
parameter signed W59TO31 = 0;
parameter signed W59TO32 = 0;
parameter signed W59TO33 = 0;
parameter signed W59TO34 = 0;
parameter signed W59TO35 = 0;
parameter signed W59TO36 = 0;
parameter signed W59TO37 = 0;
parameter signed W59TO38 = 0;
parameter signed W59TO39 = 0;
parameter signed W59TO40 = 0;
parameter signed W59TO41 = 0;
parameter signed W59TO42 = 0;
parameter signed W59TO43 = 0;
parameter signed W59TO44 = 0;
parameter signed W59TO45 = 0;
parameter signed W59TO46 = 0;
parameter signed W59TO47 = 0;
parameter signed W59TO48 = 0;
parameter signed W59TO49 = 0;
parameter signed W59TO50 = 0;
parameter signed W59TO51 = 0;
parameter signed W59TO52 = 0;
parameter signed W59TO53 = 0;
parameter signed W59TO54 = 0;
parameter signed W59TO55 = 0;
parameter signed W59TO56 = 0;
parameter signed W59TO57 = 0;
parameter signed W59TO58 = 0;
parameter signed W59TO59 = 0;
parameter signed W59TO60 = 0;
parameter signed W59TO61 = 0;
parameter signed W59TO62 = 0;
parameter signed W59TO63 = 0;
parameter signed W60TO0 = 0;
parameter signed W60TO1 = 0;
parameter signed W60TO2 = 0;
parameter signed W60TO3 = 0;
parameter signed W60TO4 = 0;
parameter signed W60TO5 = 0;
parameter signed W60TO6 = 0;
parameter signed W60TO7 = 0;
parameter signed W60TO8 = 0;
parameter signed W60TO9 = 0;
parameter signed W60TO10 = 0;
parameter signed W60TO11 = 0;
parameter signed W60TO12 = 0;
parameter signed W60TO13 = 0;
parameter signed W60TO14 = 0;
parameter signed W60TO15 = 0;
parameter signed W60TO16 = 0;
parameter signed W60TO17 = 0;
parameter signed W60TO18 = 0;
parameter signed W60TO19 = 0;
parameter signed W60TO20 = 0;
parameter signed W60TO21 = 0;
parameter signed W60TO22 = 0;
parameter signed W60TO23 = 0;
parameter signed W60TO24 = 0;
parameter signed W60TO25 = 0;
parameter signed W60TO26 = 0;
parameter signed W60TO27 = 0;
parameter signed W60TO28 = 0;
parameter signed W60TO29 = 0;
parameter signed W60TO30 = 0;
parameter signed W60TO31 = 0;
parameter signed W60TO32 = 0;
parameter signed W60TO33 = 0;
parameter signed W60TO34 = 0;
parameter signed W60TO35 = 0;
parameter signed W60TO36 = 0;
parameter signed W60TO37 = 0;
parameter signed W60TO38 = 0;
parameter signed W60TO39 = 0;
parameter signed W60TO40 = 0;
parameter signed W60TO41 = 0;
parameter signed W60TO42 = 0;
parameter signed W60TO43 = 0;
parameter signed W60TO44 = 0;
parameter signed W60TO45 = 0;
parameter signed W60TO46 = 0;
parameter signed W60TO47 = 0;
parameter signed W60TO48 = 0;
parameter signed W60TO49 = 0;
parameter signed W60TO50 = 0;
parameter signed W60TO51 = 0;
parameter signed W60TO52 = 0;
parameter signed W60TO53 = 0;
parameter signed W60TO54 = 0;
parameter signed W60TO55 = 0;
parameter signed W60TO56 = 0;
parameter signed W60TO57 = 0;
parameter signed W60TO58 = 0;
parameter signed W60TO59 = 0;
parameter signed W60TO60 = 0;
parameter signed W60TO61 = 0;
parameter signed W60TO62 = 0;
parameter signed W60TO63 = 0;
parameter signed W61TO0 = 0;
parameter signed W61TO1 = 0;
parameter signed W61TO2 = 0;
parameter signed W61TO3 = 0;
parameter signed W61TO4 = 0;
parameter signed W61TO5 = 0;
parameter signed W61TO6 = 0;
parameter signed W61TO7 = 0;
parameter signed W61TO8 = 0;
parameter signed W61TO9 = 0;
parameter signed W61TO10 = 0;
parameter signed W61TO11 = 0;
parameter signed W61TO12 = 0;
parameter signed W61TO13 = 0;
parameter signed W61TO14 = 0;
parameter signed W61TO15 = 0;
parameter signed W61TO16 = 0;
parameter signed W61TO17 = 0;
parameter signed W61TO18 = 0;
parameter signed W61TO19 = 0;
parameter signed W61TO20 = 0;
parameter signed W61TO21 = 0;
parameter signed W61TO22 = 0;
parameter signed W61TO23 = 0;
parameter signed W61TO24 = 0;
parameter signed W61TO25 = 0;
parameter signed W61TO26 = 0;
parameter signed W61TO27 = 0;
parameter signed W61TO28 = 0;
parameter signed W61TO29 = 0;
parameter signed W61TO30 = 0;
parameter signed W61TO31 = 0;
parameter signed W61TO32 = 0;
parameter signed W61TO33 = 0;
parameter signed W61TO34 = 0;
parameter signed W61TO35 = 0;
parameter signed W61TO36 = 0;
parameter signed W61TO37 = 0;
parameter signed W61TO38 = 0;
parameter signed W61TO39 = 0;
parameter signed W61TO40 = 0;
parameter signed W61TO41 = 0;
parameter signed W61TO42 = 0;
parameter signed W61TO43 = 0;
parameter signed W61TO44 = 0;
parameter signed W61TO45 = 0;
parameter signed W61TO46 = 0;
parameter signed W61TO47 = 0;
parameter signed W61TO48 = 0;
parameter signed W61TO49 = 0;
parameter signed W61TO50 = 0;
parameter signed W61TO51 = 0;
parameter signed W61TO52 = 0;
parameter signed W61TO53 = 0;
parameter signed W61TO54 = 0;
parameter signed W61TO55 = 0;
parameter signed W61TO56 = 0;
parameter signed W61TO57 = 0;
parameter signed W61TO58 = 0;
parameter signed W61TO59 = 0;
parameter signed W61TO60 = 0;
parameter signed W61TO61 = 0;
parameter signed W61TO62 = 0;
parameter signed W61TO63 = 0;
parameter signed W62TO0 = 0;
parameter signed W62TO1 = 0;
parameter signed W62TO2 = 0;
parameter signed W62TO3 = 0;
parameter signed W62TO4 = 0;
parameter signed W62TO5 = 0;
parameter signed W62TO6 = 0;
parameter signed W62TO7 = 0;
parameter signed W62TO8 = 0;
parameter signed W62TO9 = 0;
parameter signed W62TO10 = 0;
parameter signed W62TO11 = 0;
parameter signed W62TO12 = 0;
parameter signed W62TO13 = 0;
parameter signed W62TO14 = 0;
parameter signed W62TO15 = 0;
parameter signed W62TO16 = 0;
parameter signed W62TO17 = 0;
parameter signed W62TO18 = 0;
parameter signed W62TO19 = 0;
parameter signed W62TO20 = 0;
parameter signed W62TO21 = 0;
parameter signed W62TO22 = 0;
parameter signed W62TO23 = 0;
parameter signed W62TO24 = 0;
parameter signed W62TO25 = 0;
parameter signed W62TO26 = 0;
parameter signed W62TO27 = 0;
parameter signed W62TO28 = 0;
parameter signed W62TO29 = 0;
parameter signed W62TO30 = 0;
parameter signed W62TO31 = 0;
parameter signed W62TO32 = 0;
parameter signed W62TO33 = 0;
parameter signed W62TO34 = 0;
parameter signed W62TO35 = 0;
parameter signed W62TO36 = 0;
parameter signed W62TO37 = 0;
parameter signed W62TO38 = 0;
parameter signed W62TO39 = 0;
parameter signed W62TO40 = 0;
parameter signed W62TO41 = 0;
parameter signed W62TO42 = 0;
parameter signed W62TO43 = 0;
parameter signed W62TO44 = 0;
parameter signed W62TO45 = 0;
parameter signed W62TO46 = 0;
parameter signed W62TO47 = 0;
parameter signed W62TO48 = 0;
parameter signed W62TO49 = 0;
parameter signed W62TO50 = 0;
parameter signed W62TO51 = 0;
parameter signed W62TO52 = 0;
parameter signed W62TO53 = 0;
parameter signed W62TO54 = 0;
parameter signed W62TO55 = 0;
parameter signed W62TO56 = 0;
parameter signed W62TO57 = 0;
parameter signed W62TO58 = 0;
parameter signed W62TO59 = 0;
parameter signed W62TO60 = 0;
parameter signed W62TO61 = 0;
parameter signed W62TO62 = 0;
parameter signed W62TO63 = 0;
parameter signed W63TO0 = 0;
parameter signed W63TO1 = 0;
parameter signed W63TO2 = 0;
parameter signed W63TO3 = 0;
parameter signed W63TO4 = 0;
parameter signed W63TO5 = 0;
parameter signed W63TO6 = 0;
parameter signed W63TO7 = 0;
parameter signed W63TO8 = 0;
parameter signed W63TO9 = 0;
parameter signed W63TO10 = 0;
parameter signed W63TO11 = 0;
parameter signed W63TO12 = 0;
parameter signed W63TO13 = 0;
parameter signed W63TO14 = 0;
parameter signed W63TO15 = 0;
parameter signed W63TO16 = 0;
parameter signed W63TO17 = 0;
parameter signed W63TO18 = 0;
parameter signed W63TO19 = 0;
parameter signed W63TO20 = 0;
parameter signed W63TO21 = 0;
parameter signed W63TO22 = 0;
parameter signed W63TO23 = 0;
parameter signed W63TO24 = 0;
parameter signed W63TO25 = 0;
parameter signed W63TO26 = 0;
parameter signed W63TO27 = 0;
parameter signed W63TO28 = 0;
parameter signed W63TO29 = 0;
parameter signed W63TO30 = 0;
parameter signed W63TO31 = 0;
parameter signed W63TO32 = 0;
parameter signed W63TO33 = 0;
parameter signed W63TO34 = 0;
parameter signed W63TO35 = 0;
parameter signed W63TO36 = 0;
parameter signed W63TO37 = 0;
parameter signed W63TO38 = 0;
parameter signed W63TO39 = 0;
parameter signed W63TO40 = 0;
parameter signed W63TO41 = 0;
parameter signed W63TO42 = 0;
parameter signed W63TO43 = 0;
parameter signed W63TO44 = 0;
parameter signed W63TO45 = 0;
parameter signed W63TO46 = 0;
parameter signed W63TO47 = 0;
parameter signed W63TO48 = 0;
parameter signed W63TO49 = 0;
parameter signed W63TO50 = 0;
parameter signed W63TO51 = 0;
parameter signed W63TO52 = 0;
parameter signed W63TO53 = 0;
parameter signed W63TO54 = 0;
parameter signed W63TO55 = 0;
parameter signed W63TO56 = 0;
parameter signed W63TO57 = 0;
parameter signed W63TO58 = 0;
parameter signed W63TO59 = 0;
parameter signed W63TO60 = 0;
parameter signed W63TO61 = 0;
parameter signed W63TO62 = 0;
parameter signed W63TO63 = 0;
parameter signed W64TO0 = 0;
parameter signed W64TO1 = 0;
parameter signed W64TO2 = 0;
parameter signed W64TO3 = 0;
parameter signed W64TO4 = 0;
parameter signed W64TO5 = 0;
parameter signed W64TO6 = 0;
parameter signed W64TO7 = 0;
parameter signed W64TO8 = 0;
parameter signed W64TO9 = 0;
parameter signed W64TO10 = 0;
parameter signed W64TO11 = 0;
parameter signed W64TO12 = 0;
parameter signed W64TO13 = 0;
parameter signed W64TO14 = 0;
parameter signed W64TO15 = 0;
parameter signed W64TO16 = 0;
parameter signed W64TO17 = 0;
parameter signed W64TO18 = 0;
parameter signed W64TO19 = 0;
parameter signed W64TO20 = 0;
parameter signed W64TO21 = 0;
parameter signed W64TO22 = 0;
parameter signed W64TO23 = 0;
parameter signed W64TO24 = 0;
parameter signed W64TO25 = 0;
parameter signed W64TO26 = 0;
parameter signed W64TO27 = 0;
parameter signed W64TO28 = 0;
parameter signed W64TO29 = 0;
parameter signed W64TO30 = 0;
parameter signed W64TO31 = 0;
parameter signed W64TO32 = 0;
parameter signed W64TO33 = 0;
parameter signed W64TO34 = 0;
parameter signed W64TO35 = 0;
parameter signed W64TO36 = 0;
parameter signed W64TO37 = 0;
parameter signed W64TO38 = 0;
parameter signed W64TO39 = 0;
parameter signed W64TO40 = 0;
parameter signed W64TO41 = 0;
parameter signed W64TO42 = 0;
parameter signed W64TO43 = 0;
parameter signed W64TO44 = 0;
parameter signed W64TO45 = 0;
parameter signed W64TO46 = 0;
parameter signed W64TO47 = 0;
parameter signed W64TO48 = 0;
parameter signed W64TO49 = 0;
parameter signed W64TO50 = 0;
parameter signed W64TO51 = 0;
parameter signed W64TO52 = 0;
parameter signed W64TO53 = 0;
parameter signed W64TO54 = 0;
parameter signed W64TO55 = 0;
parameter signed W64TO56 = 0;
parameter signed W64TO57 = 0;
parameter signed W64TO58 = 0;
parameter signed W64TO59 = 0;
parameter signed W64TO60 = 0;
parameter signed W64TO61 = 0;
parameter signed W64TO62 = 0;
parameter signed W64TO63 = 0;

input wire clk;
input wire rst;

input signed [63:0] in0;
input signed [63:0] in1;
input signed [63:0] in2;
input signed [63:0] in3;
input signed [63:0] in4;
input signed [63:0] in5;
input signed [63:0] in6;
input signed [63:0] in7;
input signed [63:0] in8;
input signed [63:0] in9;
input signed [63:0] in10;
input signed [63:0] in11;
input signed [63:0] in12;
input signed [63:0] in13;
input signed [63:0] in14;
input signed [63:0] in15;
input signed [63:0] in16;
input signed [63:0] in17;
input signed [63:0] in18;
input signed [63:0] in19;
input signed [63:0] in20;
input signed [63:0] in21;
input signed [63:0] in22;
input signed [63:0] in23;
input signed [63:0] in24;
input signed [63:0] in25;
input signed [63:0] in26;
input signed [63:0] in27;
input signed [63:0] in28;
input signed [63:0] in29;
input signed [63:0] in30;
input signed [63:0] in31;
input signed [63:0] in32;
input signed [63:0] in33;
input signed [63:0] in34;
input signed [63:0] in35;
input signed [63:0] in36;
input signed [63:0] in37;
input signed [63:0] in38;
input signed [63:0] in39;
input signed [63:0] in40;
input signed [63:0] in41;
input signed [63:0] in42;
input signed [63:0] in43;
input signed [63:0] in44;
input signed [63:0] in45;
input signed [63:0] in46;
input signed [63:0] in47;
input signed [63:0] in48;
input signed [63:0] in49;
input signed [63:0] in50;
input signed [63:0] in51;
input signed [63:0] in52;
input signed [63:0] in53;
input signed [63:0] in54;
input signed [63:0] in55;
input signed [63:0] in56;
input signed [63:0] in57;
input signed [63:0] in58;
input signed [63:0] in59;
input signed [63:0] in60;
input signed [63:0] in61;
input signed [63:0] in62;
input signed [63:0] in63;
input signed [63:0] in64;

output signed [63:0] out0;
output signed [63:0] out1;
output signed [63:0] out2;
output signed [63:0] out3;
output signed [63:0] out4;
output signed [63:0] out5;
output signed [63:0] out6;
output signed [63:0] out7;
output signed [63:0] out8;
output signed [63:0] out9;
output signed [63:0] out10;
output signed [63:0] out11;
output signed [63:0] out12;
output signed [63:0] out13;
output signed [63:0] out14;
output signed [63:0] out15;
output signed [63:0] out16;
output signed [63:0] out17;
output signed [63:0] out18;
output signed [63:0] out19;
output signed [63:0] out20;
output signed [63:0] out21;
output signed [63:0] out22;
output signed [63:0] out23;
output signed [63:0] out24;
output signed [63:0] out25;
output signed [63:0] out26;
output signed [63:0] out27;
output signed [63:0] out28;
output signed [63:0] out29;
output signed [63:0] out30;
output signed [63:0] out31;
output signed [63:0] out32;
output signed [63:0] out33;
output signed [63:0] out34;
output signed [63:0] out35;
output signed [63:0] out36;
output signed [63:0] out37;
output signed [63:0] out38;
output signed [63:0] out39;
output signed [63:0] out40;
output signed [63:0] out41;
output signed [63:0] out42;
output signed [63:0] out43;
output signed [63:0] out44;
output signed [63:0] out45;
output signed [63:0] out46;
output signed [63:0] out47;
output signed [63:0] out48;
output signed [63:0] out49;
output signed [63:0] out50;
output signed [63:0] out51;
output signed [63:0] out52;
output signed [63:0] out53;
output signed [63:0] out54;
output signed [63:0] out55;
output signed [63:0] out56;
output signed [63:0] out57;
output signed [63:0] out58;
output signed [63:0] out59;
output signed [63:0] out60;
output signed [63:0] out61;
output signed [63:0] out62;
output signed [63:0] out63;

neuron65in #(.BIAS(BIAS0), .W0(W0TO0), .W1(W1TO0), .W2(W2TO0), .W3(W3TO0), .W4(W4TO0), .W5(W5TO0), .W6(W6TO0), .W7(W7TO0), .W8(W8TO0), .W9(W9TO0), .W10(W10TO0), .W11(W11TO0), .W12(W12TO0), .W13(W13TO0), .W14(W14TO0), .W15(W15TO0), .W16(W16TO0), .W17(W17TO0), .W18(W18TO0), .W19(W19TO0), .W20(W20TO0), .W21(W21TO0), .W22(W22TO0), .W23(W23TO0), .W24(W24TO0), .W25(W25TO0), .W26(W26TO0), .W27(W27TO0), .W28(W28TO0), .W29(W29TO0), .W30(W30TO0), .W31(W31TO0), .W32(W32TO0), .W33(W33TO0), .W34(W34TO0), .W35(W35TO0), .W36(W36TO0), .W37(W37TO0), .W38(W38TO0), .W39(W39TO0), .W40(W40TO0), .W41(W41TO0), .W42(W42TO0), .W43(W43TO0), .W44(W44TO0), .W45(W45TO0), .W46(W46TO0), .W47(W47TO0), .W48(W48TO0), .W49(W49TO0), .W50(W50TO0), .W51(W51TO0), .W52(W52TO0), .W53(W53TO0), .W54(W54TO0), .W55(W55TO0), .W56(W56TO0), .W57(W57TO0), .W58(W58TO0), .W59(W59TO0), .W60(W60TO0), .W61(W61TO0), .W62(W62TO0), .W63(W63TO0), .W64(W64TO0)) neuron0(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out0));
neuron65in #(.BIAS(BIAS1), .W0(W0TO1), .W1(W1TO1), .W2(W2TO1), .W3(W3TO1), .W4(W4TO1), .W5(W5TO1), .W6(W6TO1), .W7(W7TO1), .W8(W8TO1), .W9(W9TO1), .W10(W10TO1), .W11(W11TO1), .W12(W12TO1), .W13(W13TO1), .W14(W14TO1), .W15(W15TO1), .W16(W16TO1), .W17(W17TO1), .W18(W18TO1), .W19(W19TO1), .W20(W20TO1), .W21(W21TO1), .W22(W22TO1), .W23(W23TO1), .W24(W24TO1), .W25(W25TO1), .W26(W26TO1), .W27(W27TO1), .W28(W28TO1), .W29(W29TO1), .W30(W30TO1), .W31(W31TO1), .W32(W32TO1), .W33(W33TO1), .W34(W34TO1), .W35(W35TO1), .W36(W36TO1), .W37(W37TO1), .W38(W38TO1), .W39(W39TO1), .W40(W40TO1), .W41(W41TO1), .W42(W42TO1), .W43(W43TO1), .W44(W44TO1), .W45(W45TO1), .W46(W46TO1), .W47(W47TO1), .W48(W48TO1), .W49(W49TO1), .W50(W50TO1), .W51(W51TO1), .W52(W52TO1), .W53(W53TO1), .W54(W54TO1), .W55(W55TO1), .W56(W56TO1), .W57(W57TO1), .W58(W58TO1), .W59(W59TO1), .W60(W60TO1), .W61(W61TO1), .W62(W62TO1), .W63(W63TO1), .W64(W64TO1)) neuron1(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out1));
neuron65in #(.BIAS(BIAS2), .W0(W0TO2), .W1(W1TO2), .W2(W2TO2), .W3(W3TO2), .W4(W4TO2), .W5(W5TO2), .W6(W6TO2), .W7(W7TO2), .W8(W8TO2), .W9(W9TO2), .W10(W10TO2), .W11(W11TO2), .W12(W12TO2), .W13(W13TO2), .W14(W14TO2), .W15(W15TO2), .W16(W16TO2), .W17(W17TO2), .W18(W18TO2), .W19(W19TO2), .W20(W20TO2), .W21(W21TO2), .W22(W22TO2), .W23(W23TO2), .W24(W24TO2), .W25(W25TO2), .W26(W26TO2), .W27(W27TO2), .W28(W28TO2), .W29(W29TO2), .W30(W30TO2), .W31(W31TO2), .W32(W32TO2), .W33(W33TO2), .W34(W34TO2), .W35(W35TO2), .W36(W36TO2), .W37(W37TO2), .W38(W38TO2), .W39(W39TO2), .W40(W40TO2), .W41(W41TO2), .W42(W42TO2), .W43(W43TO2), .W44(W44TO2), .W45(W45TO2), .W46(W46TO2), .W47(W47TO2), .W48(W48TO2), .W49(W49TO2), .W50(W50TO2), .W51(W51TO2), .W52(W52TO2), .W53(W53TO2), .W54(W54TO2), .W55(W55TO2), .W56(W56TO2), .W57(W57TO2), .W58(W58TO2), .W59(W59TO2), .W60(W60TO2), .W61(W61TO2), .W62(W62TO2), .W63(W63TO2), .W64(W64TO2)) neuron2(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out2));
neuron65in #(.BIAS(BIAS3), .W0(W0TO3), .W1(W1TO3), .W2(W2TO3), .W3(W3TO3), .W4(W4TO3), .W5(W5TO3), .W6(W6TO3), .W7(W7TO3), .W8(W8TO3), .W9(W9TO3), .W10(W10TO3), .W11(W11TO3), .W12(W12TO3), .W13(W13TO3), .W14(W14TO3), .W15(W15TO3), .W16(W16TO3), .W17(W17TO3), .W18(W18TO3), .W19(W19TO3), .W20(W20TO3), .W21(W21TO3), .W22(W22TO3), .W23(W23TO3), .W24(W24TO3), .W25(W25TO3), .W26(W26TO3), .W27(W27TO3), .W28(W28TO3), .W29(W29TO3), .W30(W30TO3), .W31(W31TO3), .W32(W32TO3), .W33(W33TO3), .W34(W34TO3), .W35(W35TO3), .W36(W36TO3), .W37(W37TO3), .W38(W38TO3), .W39(W39TO3), .W40(W40TO3), .W41(W41TO3), .W42(W42TO3), .W43(W43TO3), .W44(W44TO3), .W45(W45TO3), .W46(W46TO3), .W47(W47TO3), .W48(W48TO3), .W49(W49TO3), .W50(W50TO3), .W51(W51TO3), .W52(W52TO3), .W53(W53TO3), .W54(W54TO3), .W55(W55TO3), .W56(W56TO3), .W57(W57TO3), .W58(W58TO3), .W59(W59TO3), .W60(W60TO3), .W61(W61TO3), .W62(W62TO3), .W63(W63TO3), .W64(W64TO3)) neuron3(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out3));
neuron65in #(.BIAS(BIAS4), .W0(W0TO4), .W1(W1TO4), .W2(W2TO4), .W3(W3TO4), .W4(W4TO4), .W5(W5TO4), .W6(W6TO4), .W7(W7TO4), .W8(W8TO4), .W9(W9TO4), .W10(W10TO4), .W11(W11TO4), .W12(W12TO4), .W13(W13TO4), .W14(W14TO4), .W15(W15TO4), .W16(W16TO4), .W17(W17TO4), .W18(W18TO4), .W19(W19TO4), .W20(W20TO4), .W21(W21TO4), .W22(W22TO4), .W23(W23TO4), .W24(W24TO4), .W25(W25TO4), .W26(W26TO4), .W27(W27TO4), .W28(W28TO4), .W29(W29TO4), .W30(W30TO4), .W31(W31TO4), .W32(W32TO4), .W33(W33TO4), .W34(W34TO4), .W35(W35TO4), .W36(W36TO4), .W37(W37TO4), .W38(W38TO4), .W39(W39TO4), .W40(W40TO4), .W41(W41TO4), .W42(W42TO4), .W43(W43TO4), .W44(W44TO4), .W45(W45TO4), .W46(W46TO4), .W47(W47TO4), .W48(W48TO4), .W49(W49TO4), .W50(W50TO4), .W51(W51TO4), .W52(W52TO4), .W53(W53TO4), .W54(W54TO4), .W55(W55TO4), .W56(W56TO4), .W57(W57TO4), .W58(W58TO4), .W59(W59TO4), .W60(W60TO4), .W61(W61TO4), .W62(W62TO4), .W63(W63TO4), .W64(W64TO4)) neuron4(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out4));
neuron65in #(.BIAS(BIAS5), .W0(W0TO5), .W1(W1TO5), .W2(W2TO5), .W3(W3TO5), .W4(W4TO5), .W5(W5TO5), .W6(W6TO5), .W7(W7TO5), .W8(W8TO5), .W9(W9TO5), .W10(W10TO5), .W11(W11TO5), .W12(W12TO5), .W13(W13TO5), .W14(W14TO5), .W15(W15TO5), .W16(W16TO5), .W17(W17TO5), .W18(W18TO5), .W19(W19TO5), .W20(W20TO5), .W21(W21TO5), .W22(W22TO5), .W23(W23TO5), .W24(W24TO5), .W25(W25TO5), .W26(W26TO5), .W27(W27TO5), .W28(W28TO5), .W29(W29TO5), .W30(W30TO5), .W31(W31TO5), .W32(W32TO5), .W33(W33TO5), .W34(W34TO5), .W35(W35TO5), .W36(W36TO5), .W37(W37TO5), .W38(W38TO5), .W39(W39TO5), .W40(W40TO5), .W41(W41TO5), .W42(W42TO5), .W43(W43TO5), .W44(W44TO5), .W45(W45TO5), .W46(W46TO5), .W47(W47TO5), .W48(W48TO5), .W49(W49TO5), .W50(W50TO5), .W51(W51TO5), .W52(W52TO5), .W53(W53TO5), .W54(W54TO5), .W55(W55TO5), .W56(W56TO5), .W57(W57TO5), .W58(W58TO5), .W59(W59TO5), .W60(W60TO5), .W61(W61TO5), .W62(W62TO5), .W63(W63TO5), .W64(W64TO5)) neuron5(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out5));
neuron65in #(.BIAS(BIAS6), .W0(W0TO6), .W1(W1TO6), .W2(W2TO6), .W3(W3TO6), .W4(W4TO6), .W5(W5TO6), .W6(W6TO6), .W7(W7TO6), .W8(W8TO6), .W9(W9TO6), .W10(W10TO6), .W11(W11TO6), .W12(W12TO6), .W13(W13TO6), .W14(W14TO6), .W15(W15TO6), .W16(W16TO6), .W17(W17TO6), .W18(W18TO6), .W19(W19TO6), .W20(W20TO6), .W21(W21TO6), .W22(W22TO6), .W23(W23TO6), .W24(W24TO6), .W25(W25TO6), .W26(W26TO6), .W27(W27TO6), .W28(W28TO6), .W29(W29TO6), .W30(W30TO6), .W31(W31TO6), .W32(W32TO6), .W33(W33TO6), .W34(W34TO6), .W35(W35TO6), .W36(W36TO6), .W37(W37TO6), .W38(W38TO6), .W39(W39TO6), .W40(W40TO6), .W41(W41TO6), .W42(W42TO6), .W43(W43TO6), .W44(W44TO6), .W45(W45TO6), .W46(W46TO6), .W47(W47TO6), .W48(W48TO6), .W49(W49TO6), .W50(W50TO6), .W51(W51TO6), .W52(W52TO6), .W53(W53TO6), .W54(W54TO6), .W55(W55TO6), .W56(W56TO6), .W57(W57TO6), .W58(W58TO6), .W59(W59TO6), .W60(W60TO6), .W61(W61TO6), .W62(W62TO6), .W63(W63TO6), .W64(W64TO6)) neuron6(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out6));
neuron65in #(.BIAS(BIAS7), .W0(W0TO7), .W1(W1TO7), .W2(W2TO7), .W3(W3TO7), .W4(W4TO7), .W5(W5TO7), .W6(W6TO7), .W7(W7TO7), .W8(W8TO7), .W9(W9TO7), .W10(W10TO7), .W11(W11TO7), .W12(W12TO7), .W13(W13TO7), .W14(W14TO7), .W15(W15TO7), .W16(W16TO7), .W17(W17TO7), .W18(W18TO7), .W19(W19TO7), .W20(W20TO7), .W21(W21TO7), .W22(W22TO7), .W23(W23TO7), .W24(W24TO7), .W25(W25TO7), .W26(W26TO7), .W27(W27TO7), .W28(W28TO7), .W29(W29TO7), .W30(W30TO7), .W31(W31TO7), .W32(W32TO7), .W33(W33TO7), .W34(W34TO7), .W35(W35TO7), .W36(W36TO7), .W37(W37TO7), .W38(W38TO7), .W39(W39TO7), .W40(W40TO7), .W41(W41TO7), .W42(W42TO7), .W43(W43TO7), .W44(W44TO7), .W45(W45TO7), .W46(W46TO7), .W47(W47TO7), .W48(W48TO7), .W49(W49TO7), .W50(W50TO7), .W51(W51TO7), .W52(W52TO7), .W53(W53TO7), .W54(W54TO7), .W55(W55TO7), .W56(W56TO7), .W57(W57TO7), .W58(W58TO7), .W59(W59TO7), .W60(W60TO7), .W61(W61TO7), .W62(W62TO7), .W63(W63TO7), .W64(W64TO7)) neuron7(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out7));
neuron65in #(.BIAS(BIAS8), .W0(W0TO8), .W1(W1TO8), .W2(W2TO8), .W3(W3TO8), .W4(W4TO8), .W5(W5TO8), .W6(W6TO8), .W7(W7TO8), .W8(W8TO8), .W9(W9TO8), .W10(W10TO8), .W11(W11TO8), .W12(W12TO8), .W13(W13TO8), .W14(W14TO8), .W15(W15TO8), .W16(W16TO8), .W17(W17TO8), .W18(W18TO8), .W19(W19TO8), .W20(W20TO8), .W21(W21TO8), .W22(W22TO8), .W23(W23TO8), .W24(W24TO8), .W25(W25TO8), .W26(W26TO8), .W27(W27TO8), .W28(W28TO8), .W29(W29TO8), .W30(W30TO8), .W31(W31TO8), .W32(W32TO8), .W33(W33TO8), .W34(W34TO8), .W35(W35TO8), .W36(W36TO8), .W37(W37TO8), .W38(W38TO8), .W39(W39TO8), .W40(W40TO8), .W41(W41TO8), .W42(W42TO8), .W43(W43TO8), .W44(W44TO8), .W45(W45TO8), .W46(W46TO8), .W47(W47TO8), .W48(W48TO8), .W49(W49TO8), .W50(W50TO8), .W51(W51TO8), .W52(W52TO8), .W53(W53TO8), .W54(W54TO8), .W55(W55TO8), .W56(W56TO8), .W57(W57TO8), .W58(W58TO8), .W59(W59TO8), .W60(W60TO8), .W61(W61TO8), .W62(W62TO8), .W63(W63TO8), .W64(W64TO8)) neuron8(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out8));
neuron65in #(.BIAS(BIAS9), .W0(W0TO9), .W1(W1TO9), .W2(W2TO9), .W3(W3TO9), .W4(W4TO9), .W5(W5TO9), .W6(W6TO9), .W7(W7TO9), .W8(W8TO9), .W9(W9TO9), .W10(W10TO9), .W11(W11TO9), .W12(W12TO9), .W13(W13TO9), .W14(W14TO9), .W15(W15TO9), .W16(W16TO9), .W17(W17TO9), .W18(W18TO9), .W19(W19TO9), .W20(W20TO9), .W21(W21TO9), .W22(W22TO9), .W23(W23TO9), .W24(W24TO9), .W25(W25TO9), .W26(W26TO9), .W27(W27TO9), .W28(W28TO9), .W29(W29TO9), .W30(W30TO9), .W31(W31TO9), .W32(W32TO9), .W33(W33TO9), .W34(W34TO9), .W35(W35TO9), .W36(W36TO9), .W37(W37TO9), .W38(W38TO9), .W39(W39TO9), .W40(W40TO9), .W41(W41TO9), .W42(W42TO9), .W43(W43TO9), .W44(W44TO9), .W45(W45TO9), .W46(W46TO9), .W47(W47TO9), .W48(W48TO9), .W49(W49TO9), .W50(W50TO9), .W51(W51TO9), .W52(W52TO9), .W53(W53TO9), .W54(W54TO9), .W55(W55TO9), .W56(W56TO9), .W57(W57TO9), .W58(W58TO9), .W59(W59TO9), .W60(W60TO9), .W61(W61TO9), .W62(W62TO9), .W63(W63TO9), .W64(W64TO9)) neuron9(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out9));
neuron65in #(.BIAS(BIAS10), .W0(W0TO10), .W1(W1TO10), .W2(W2TO10), .W3(W3TO10), .W4(W4TO10), .W5(W5TO10), .W6(W6TO10), .W7(W7TO10), .W8(W8TO10), .W9(W9TO10), .W10(W10TO10), .W11(W11TO10), .W12(W12TO10), .W13(W13TO10), .W14(W14TO10), .W15(W15TO10), .W16(W16TO10), .W17(W17TO10), .W18(W18TO10), .W19(W19TO10), .W20(W20TO10), .W21(W21TO10), .W22(W22TO10), .W23(W23TO10), .W24(W24TO10), .W25(W25TO10), .W26(W26TO10), .W27(W27TO10), .W28(W28TO10), .W29(W29TO10), .W30(W30TO10), .W31(W31TO10), .W32(W32TO10), .W33(W33TO10), .W34(W34TO10), .W35(W35TO10), .W36(W36TO10), .W37(W37TO10), .W38(W38TO10), .W39(W39TO10), .W40(W40TO10), .W41(W41TO10), .W42(W42TO10), .W43(W43TO10), .W44(W44TO10), .W45(W45TO10), .W46(W46TO10), .W47(W47TO10), .W48(W48TO10), .W49(W49TO10), .W50(W50TO10), .W51(W51TO10), .W52(W52TO10), .W53(W53TO10), .W54(W54TO10), .W55(W55TO10), .W56(W56TO10), .W57(W57TO10), .W58(W58TO10), .W59(W59TO10), .W60(W60TO10), .W61(W61TO10), .W62(W62TO10), .W63(W63TO10), .W64(W64TO10)) neuron10(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out10));
neuron65in #(.BIAS(BIAS11), .W0(W0TO11), .W1(W1TO11), .W2(W2TO11), .W3(W3TO11), .W4(W4TO11), .W5(W5TO11), .W6(W6TO11), .W7(W7TO11), .W8(W8TO11), .W9(W9TO11), .W10(W10TO11), .W11(W11TO11), .W12(W12TO11), .W13(W13TO11), .W14(W14TO11), .W15(W15TO11), .W16(W16TO11), .W17(W17TO11), .W18(W18TO11), .W19(W19TO11), .W20(W20TO11), .W21(W21TO11), .W22(W22TO11), .W23(W23TO11), .W24(W24TO11), .W25(W25TO11), .W26(W26TO11), .W27(W27TO11), .W28(W28TO11), .W29(W29TO11), .W30(W30TO11), .W31(W31TO11), .W32(W32TO11), .W33(W33TO11), .W34(W34TO11), .W35(W35TO11), .W36(W36TO11), .W37(W37TO11), .W38(W38TO11), .W39(W39TO11), .W40(W40TO11), .W41(W41TO11), .W42(W42TO11), .W43(W43TO11), .W44(W44TO11), .W45(W45TO11), .W46(W46TO11), .W47(W47TO11), .W48(W48TO11), .W49(W49TO11), .W50(W50TO11), .W51(W51TO11), .W52(W52TO11), .W53(W53TO11), .W54(W54TO11), .W55(W55TO11), .W56(W56TO11), .W57(W57TO11), .W58(W58TO11), .W59(W59TO11), .W60(W60TO11), .W61(W61TO11), .W62(W62TO11), .W63(W63TO11), .W64(W64TO11)) neuron11(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out11));
neuron65in #(.BIAS(BIAS12), .W0(W0TO12), .W1(W1TO12), .W2(W2TO12), .W3(W3TO12), .W4(W4TO12), .W5(W5TO12), .W6(W6TO12), .W7(W7TO12), .W8(W8TO12), .W9(W9TO12), .W10(W10TO12), .W11(W11TO12), .W12(W12TO12), .W13(W13TO12), .W14(W14TO12), .W15(W15TO12), .W16(W16TO12), .W17(W17TO12), .W18(W18TO12), .W19(W19TO12), .W20(W20TO12), .W21(W21TO12), .W22(W22TO12), .W23(W23TO12), .W24(W24TO12), .W25(W25TO12), .W26(W26TO12), .W27(W27TO12), .W28(W28TO12), .W29(W29TO12), .W30(W30TO12), .W31(W31TO12), .W32(W32TO12), .W33(W33TO12), .W34(W34TO12), .W35(W35TO12), .W36(W36TO12), .W37(W37TO12), .W38(W38TO12), .W39(W39TO12), .W40(W40TO12), .W41(W41TO12), .W42(W42TO12), .W43(W43TO12), .W44(W44TO12), .W45(W45TO12), .W46(W46TO12), .W47(W47TO12), .W48(W48TO12), .W49(W49TO12), .W50(W50TO12), .W51(W51TO12), .W52(W52TO12), .W53(W53TO12), .W54(W54TO12), .W55(W55TO12), .W56(W56TO12), .W57(W57TO12), .W58(W58TO12), .W59(W59TO12), .W60(W60TO12), .W61(W61TO12), .W62(W62TO12), .W63(W63TO12), .W64(W64TO12)) neuron12(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out12));
neuron65in #(.BIAS(BIAS13), .W0(W0TO13), .W1(W1TO13), .W2(W2TO13), .W3(W3TO13), .W4(W4TO13), .W5(W5TO13), .W6(W6TO13), .W7(W7TO13), .W8(W8TO13), .W9(W9TO13), .W10(W10TO13), .W11(W11TO13), .W12(W12TO13), .W13(W13TO13), .W14(W14TO13), .W15(W15TO13), .W16(W16TO13), .W17(W17TO13), .W18(W18TO13), .W19(W19TO13), .W20(W20TO13), .W21(W21TO13), .W22(W22TO13), .W23(W23TO13), .W24(W24TO13), .W25(W25TO13), .W26(W26TO13), .W27(W27TO13), .W28(W28TO13), .W29(W29TO13), .W30(W30TO13), .W31(W31TO13), .W32(W32TO13), .W33(W33TO13), .W34(W34TO13), .W35(W35TO13), .W36(W36TO13), .W37(W37TO13), .W38(W38TO13), .W39(W39TO13), .W40(W40TO13), .W41(W41TO13), .W42(W42TO13), .W43(W43TO13), .W44(W44TO13), .W45(W45TO13), .W46(W46TO13), .W47(W47TO13), .W48(W48TO13), .W49(W49TO13), .W50(W50TO13), .W51(W51TO13), .W52(W52TO13), .W53(W53TO13), .W54(W54TO13), .W55(W55TO13), .W56(W56TO13), .W57(W57TO13), .W58(W58TO13), .W59(W59TO13), .W60(W60TO13), .W61(W61TO13), .W62(W62TO13), .W63(W63TO13), .W64(W64TO13)) neuron13(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out13));
neuron65in #(.BIAS(BIAS14), .W0(W0TO14), .W1(W1TO14), .W2(W2TO14), .W3(W3TO14), .W4(W4TO14), .W5(W5TO14), .W6(W6TO14), .W7(W7TO14), .W8(W8TO14), .W9(W9TO14), .W10(W10TO14), .W11(W11TO14), .W12(W12TO14), .W13(W13TO14), .W14(W14TO14), .W15(W15TO14), .W16(W16TO14), .W17(W17TO14), .W18(W18TO14), .W19(W19TO14), .W20(W20TO14), .W21(W21TO14), .W22(W22TO14), .W23(W23TO14), .W24(W24TO14), .W25(W25TO14), .W26(W26TO14), .W27(W27TO14), .W28(W28TO14), .W29(W29TO14), .W30(W30TO14), .W31(W31TO14), .W32(W32TO14), .W33(W33TO14), .W34(W34TO14), .W35(W35TO14), .W36(W36TO14), .W37(W37TO14), .W38(W38TO14), .W39(W39TO14), .W40(W40TO14), .W41(W41TO14), .W42(W42TO14), .W43(W43TO14), .W44(W44TO14), .W45(W45TO14), .W46(W46TO14), .W47(W47TO14), .W48(W48TO14), .W49(W49TO14), .W50(W50TO14), .W51(W51TO14), .W52(W52TO14), .W53(W53TO14), .W54(W54TO14), .W55(W55TO14), .W56(W56TO14), .W57(W57TO14), .W58(W58TO14), .W59(W59TO14), .W60(W60TO14), .W61(W61TO14), .W62(W62TO14), .W63(W63TO14), .W64(W64TO14)) neuron14(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out14));
neuron65in #(.BIAS(BIAS15), .W0(W0TO15), .W1(W1TO15), .W2(W2TO15), .W3(W3TO15), .W4(W4TO15), .W5(W5TO15), .W6(W6TO15), .W7(W7TO15), .W8(W8TO15), .W9(W9TO15), .W10(W10TO15), .W11(W11TO15), .W12(W12TO15), .W13(W13TO15), .W14(W14TO15), .W15(W15TO15), .W16(W16TO15), .W17(W17TO15), .W18(W18TO15), .W19(W19TO15), .W20(W20TO15), .W21(W21TO15), .W22(W22TO15), .W23(W23TO15), .W24(W24TO15), .W25(W25TO15), .W26(W26TO15), .W27(W27TO15), .W28(W28TO15), .W29(W29TO15), .W30(W30TO15), .W31(W31TO15), .W32(W32TO15), .W33(W33TO15), .W34(W34TO15), .W35(W35TO15), .W36(W36TO15), .W37(W37TO15), .W38(W38TO15), .W39(W39TO15), .W40(W40TO15), .W41(W41TO15), .W42(W42TO15), .W43(W43TO15), .W44(W44TO15), .W45(W45TO15), .W46(W46TO15), .W47(W47TO15), .W48(W48TO15), .W49(W49TO15), .W50(W50TO15), .W51(W51TO15), .W52(W52TO15), .W53(W53TO15), .W54(W54TO15), .W55(W55TO15), .W56(W56TO15), .W57(W57TO15), .W58(W58TO15), .W59(W59TO15), .W60(W60TO15), .W61(W61TO15), .W62(W62TO15), .W63(W63TO15), .W64(W64TO15)) neuron15(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out15));
neuron65in #(.BIAS(BIAS16), .W0(W0TO16), .W1(W1TO16), .W2(W2TO16), .W3(W3TO16), .W4(W4TO16), .W5(W5TO16), .W6(W6TO16), .W7(W7TO16), .W8(W8TO16), .W9(W9TO16), .W10(W10TO16), .W11(W11TO16), .W12(W12TO16), .W13(W13TO16), .W14(W14TO16), .W15(W15TO16), .W16(W16TO16), .W17(W17TO16), .W18(W18TO16), .W19(W19TO16), .W20(W20TO16), .W21(W21TO16), .W22(W22TO16), .W23(W23TO16), .W24(W24TO16), .W25(W25TO16), .W26(W26TO16), .W27(W27TO16), .W28(W28TO16), .W29(W29TO16), .W30(W30TO16), .W31(W31TO16), .W32(W32TO16), .W33(W33TO16), .W34(W34TO16), .W35(W35TO16), .W36(W36TO16), .W37(W37TO16), .W38(W38TO16), .W39(W39TO16), .W40(W40TO16), .W41(W41TO16), .W42(W42TO16), .W43(W43TO16), .W44(W44TO16), .W45(W45TO16), .W46(W46TO16), .W47(W47TO16), .W48(W48TO16), .W49(W49TO16), .W50(W50TO16), .W51(W51TO16), .W52(W52TO16), .W53(W53TO16), .W54(W54TO16), .W55(W55TO16), .W56(W56TO16), .W57(W57TO16), .W58(W58TO16), .W59(W59TO16), .W60(W60TO16), .W61(W61TO16), .W62(W62TO16), .W63(W63TO16), .W64(W64TO16)) neuron16(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out16));
neuron65in #(.BIAS(BIAS17), .W0(W0TO17), .W1(W1TO17), .W2(W2TO17), .W3(W3TO17), .W4(W4TO17), .W5(W5TO17), .W6(W6TO17), .W7(W7TO17), .W8(W8TO17), .W9(W9TO17), .W10(W10TO17), .W11(W11TO17), .W12(W12TO17), .W13(W13TO17), .W14(W14TO17), .W15(W15TO17), .W16(W16TO17), .W17(W17TO17), .W18(W18TO17), .W19(W19TO17), .W20(W20TO17), .W21(W21TO17), .W22(W22TO17), .W23(W23TO17), .W24(W24TO17), .W25(W25TO17), .W26(W26TO17), .W27(W27TO17), .W28(W28TO17), .W29(W29TO17), .W30(W30TO17), .W31(W31TO17), .W32(W32TO17), .W33(W33TO17), .W34(W34TO17), .W35(W35TO17), .W36(W36TO17), .W37(W37TO17), .W38(W38TO17), .W39(W39TO17), .W40(W40TO17), .W41(W41TO17), .W42(W42TO17), .W43(W43TO17), .W44(W44TO17), .W45(W45TO17), .W46(W46TO17), .W47(W47TO17), .W48(W48TO17), .W49(W49TO17), .W50(W50TO17), .W51(W51TO17), .W52(W52TO17), .W53(W53TO17), .W54(W54TO17), .W55(W55TO17), .W56(W56TO17), .W57(W57TO17), .W58(W58TO17), .W59(W59TO17), .W60(W60TO17), .W61(W61TO17), .W62(W62TO17), .W63(W63TO17), .W64(W64TO17)) neuron17(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out17));
neuron65in #(.BIAS(BIAS18), .W0(W0TO18), .W1(W1TO18), .W2(W2TO18), .W3(W3TO18), .W4(W4TO18), .W5(W5TO18), .W6(W6TO18), .W7(W7TO18), .W8(W8TO18), .W9(W9TO18), .W10(W10TO18), .W11(W11TO18), .W12(W12TO18), .W13(W13TO18), .W14(W14TO18), .W15(W15TO18), .W16(W16TO18), .W17(W17TO18), .W18(W18TO18), .W19(W19TO18), .W20(W20TO18), .W21(W21TO18), .W22(W22TO18), .W23(W23TO18), .W24(W24TO18), .W25(W25TO18), .W26(W26TO18), .W27(W27TO18), .W28(W28TO18), .W29(W29TO18), .W30(W30TO18), .W31(W31TO18), .W32(W32TO18), .W33(W33TO18), .W34(W34TO18), .W35(W35TO18), .W36(W36TO18), .W37(W37TO18), .W38(W38TO18), .W39(W39TO18), .W40(W40TO18), .W41(W41TO18), .W42(W42TO18), .W43(W43TO18), .W44(W44TO18), .W45(W45TO18), .W46(W46TO18), .W47(W47TO18), .W48(W48TO18), .W49(W49TO18), .W50(W50TO18), .W51(W51TO18), .W52(W52TO18), .W53(W53TO18), .W54(W54TO18), .W55(W55TO18), .W56(W56TO18), .W57(W57TO18), .W58(W58TO18), .W59(W59TO18), .W60(W60TO18), .W61(W61TO18), .W62(W62TO18), .W63(W63TO18), .W64(W64TO18)) neuron18(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out18));
neuron65in #(.BIAS(BIAS19), .W0(W0TO19), .W1(W1TO19), .W2(W2TO19), .W3(W3TO19), .W4(W4TO19), .W5(W5TO19), .W6(W6TO19), .W7(W7TO19), .W8(W8TO19), .W9(W9TO19), .W10(W10TO19), .W11(W11TO19), .W12(W12TO19), .W13(W13TO19), .W14(W14TO19), .W15(W15TO19), .W16(W16TO19), .W17(W17TO19), .W18(W18TO19), .W19(W19TO19), .W20(W20TO19), .W21(W21TO19), .W22(W22TO19), .W23(W23TO19), .W24(W24TO19), .W25(W25TO19), .W26(W26TO19), .W27(W27TO19), .W28(W28TO19), .W29(W29TO19), .W30(W30TO19), .W31(W31TO19), .W32(W32TO19), .W33(W33TO19), .W34(W34TO19), .W35(W35TO19), .W36(W36TO19), .W37(W37TO19), .W38(W38TO19), .W39(W39TO19), .W40(W40TO19), .W41(W41TO19), .W42(W42TO19), .W43(W43TO19), .W44(W44TO19), .W45(W45TO19), .W46(W46TO19), .W47(W47TO19), .W48(W48TO19), .W49(W49TO19), .W50(W50TO19), .W51(W51TO19), .W52(W52TO19), .W53(W53TO19), .W54(W54TO19), .W55(W55TO19), .W56(W56TO19), .W57(W57TO19), .W58(W58TO19), .W59(W59TO19), .W60(W60TO19), .W61(W61TO19), .W62(W62TO19), .W63(W63TO19), .W64(W64TO19)) neuron19(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out19));
neuron65in #(.BIAS(BIAS20), .W0(W0TO20), .W1(W1TO20), .W2(W2TO20), .W3(W3TO20), .W4(W4TO20), .W5(W5TO20), .W6(W6TO20), .W7(W7TO20), .W8(W8TO20), .W9(W9TO20), .W10(W10TO20), .W11(W11TO20), .W12(W12TO20), .W13(W13TO20), .W14(W14TO20), .W15(W15TO20), .W16(W16TO20), .W17(W17TO20), .W18(W18TO20), .W19(W19TO20), .W20(W20TO20), .W21(W21TO20), .W22(W22TO20), .W23(W23TO20), .W24(W24TO20), .W25(W25TO20), .W26(W26TO20), .W27(W27TO20), .W28(W28TO20), .W29(W29TO20), .W30(W30TO20), .W31(W31TO20), .W32(W32TO20), .W33(W33TO20), .W34(W34TO20), .W35(W35TO20), .W36(W36TO20), .W37(W37TO20), .W38(W38TO20), .W39(W39TO20), .W40(W40TO20), .W41(W41TO20), .W42(W42TO20), .W43(W43TO20), .W44(W44TO20), .W45(W45TO20), .W46(W46TO20), .W47(W47TO20), .W48(W48TO20), .W49(W49TO20), .W50(W50TO20), .W51(W51TO20), .W52(W52TO20), .W53(W53TO20), .W54(W54TO20), .W55(W55TO20), .W56(W56TO20), .W57(W57TO20), .W58(W58TO20), .W59(W59TO20), .W60(W60TO20), .W61(W61TO20), .W62(W62TO20), .W63(W63TO20), .W64(W64TO20)) neuron20(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out20));
neuron65in #(.BIAS(BIAS21), .W0(W0TO21), .W1(W1TO21), .W2(W2TO21), .W3(W3TO21), .W4(W4TO21), .W5(W5TO21), .W6(W6TO21), .W7(W7TO21), .W8(W8TO21), .W9(W9TO21), .W10(W10TO21), .W11(W11TO21), .W12(W12TO21), .W13(W13TO21), .W14(W14TO21), .W15(W15TO21), .W16(W16TO21), .W17(W17TO21), .W18(W18TO21), .W19(W19TO21), .W20(W20TO21), .W21(W21TO21), .W22(W22TO21), .W23(W23TO21), .W24(W24TO21), .W25(W25TO21), .W26(W26TO21), .W27(W27TO21), .W28(W28TO21), .W29(W29TO21), .W30(W30TO21), .W31(W31TO21), .W32(W32TO21), .W33(W33TO21), .W34(W34TO21), .W35(W35TO21), .W36(W36TO21), .W37(W37TO21), .W38(W38TO21), .W39(W39TO21), .W40(W40TO21), .W41(W41TO21), .W42(W42TO21), .W43(W43TO21), .W44(W44TO21), .W45(W45TO21), .W46(W46TO21), .W47(W47TO21), .W48(W48TO21), .W49(W49TO21), .W50(W50TO21), .W51(W51TO21), .W52(W52TO21), .W53(W53TO21), .W54(W54TO21), .W55(W55TO21), .W56(W56TO21), .W57(W57TO21), .W58(W58TO21), .W59(W59TO21), .W60(W60TO21), .W61(W61TO21), .W62(W62TO21), .W63(W63TO21), .W64(W64TO21)) neuron21(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out21));
neuron65in #(.BIAS(BIAS22), .W0(W0TO22), .W1(W1TO22), .W2(W2TO22), .W3(W3TO22), .W4(W4TO22), .W5(W5TO22), .W6(W6TO22), .W7(W7TO22), .W8(W8TO22), .W9(W9TO22), .W10(W10TO22), .W11(W11TO22), .W12(W12TO22), .W13(W13TO22), .W14(W14TO22), .W15(W15TO22), .W16(W16TO22), .W17(W17TO22), .W18(W18TO22), .W19(W19TO22), .W20(W20TO22), .W21(W21TO22), .W22(W22TO22), .W23(W23TO22), .W24(W24TO22), .W25(W25TO22), .W26(W26TO22), .W27(W27TO22), .W28(W28TO22), .W29(W29TO22), .W30(W30TO22), .W31(W31TO22), .W32(W32TO22), .W33(W33TO22), .W34(W34TO22), .W35(W35TO22), .W36(W36TO22), .W37(W37TO22), .W38(W38TO22), .W39(W39TO22), .W40(W40TO22), .W41(W41TO22), .W42(W42TO22), .W43(W43TO22), .W44(W44TO22), .W45(W45TO22), .W46(W46TO22), .W47(W47TO22), .W48(W48TO22), .W49(W49TO22), .W50(W50TO22), .W51(W51TO22), .W52(W52TO22), .W53(W53TO22), .W54(W54TO22), .W55(W55TO22), .W56(W56TO22), .W57(W57TO22), .W58(W58TO22), .W59(W59TO22), .W60(W60TO22), .W61(W61TO22), .W62(W62TO22), .W63(W63TO22), .W64(W64TO22)) neuron22(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out22));
neuron65in #(.BIAS(BIAS23), .W0(W0TO23), .W1(W1TO23), .W2(W2TO23), .W3(W3TO23), .W4(W4TO23), .W5(W5TO23), .W6(W6TO23), .W7(W7TO23), .W8(W8TO23), .W9(W9TO23), .W10(W10TO23), .W11(W11TO23), .W12(W12TO23), .W13(W13TO23), .W14(W14TO23), .W15(W15TO23), .W16(W16TO23), .W17(W17TO23), .W18(W18TO23), .W19(W19TO23), .W20(W20TO23), .W21(W21TO23), .W22(W22TO23), .W23(W23TO23), .W24(W24TO23), .W25(W25TO23), .W26(W26TO23), .W27(W27TO23), .W28(W28TO23), .W29(W29TO23), .W30(W30TO23), .W31(W31TO23), .W32(W32TO23), .W33(W33TO23), .W34(W34TO23), .W35(W35TO23), .W36(W36TO23), .W37(W37TO23), .W38(W38TO23), .W39(W39TO23), .W40(W40TO23), .W41(W41TO23), .W42(W42TO23), .W43(W43TO23), .W44(W44TO23), .W45(W45TO23), .W46(W46TO23), .W47(W47TO23), .W48(W48TO23), .W49(W49TO23), .W50(W50TO23), .W51(W51TO23), .W52(W52TO23), .W53(W53TO23), .W54(W54TO23), .W55(W55TO23), .W56(W56TO23), .W57(W57TO23), .W58(W58TO23), .W59(W59TO23), .W60(W60TO23), .W61(W61TO23), .W62(W62TO23), .W63(W63TO23), .W64(W64TO23)) neuron23(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out23));
neuron65in #(.BIAS(BIAS24), .W0(W0TO24), .W1(W1TO24), .W2(W2TO24), .W3(W3TO24), .W4(W4TO24), .W5(W5TO24), .W6(W6TO24), .W7(W7TO24), .W8(W8TO24), .W9(W9TO24), .W10(W10TO24), .W11(W11TO24), .W12(W12TO24), .W13(W13TO24), .W14(W14TO24), .W15(W15TO24), .W16(W16TO24), .W17(W17TO24), .W18(W18TO24), .W19(W19TO24), .W20(W20TO24), .W21(W21TO24), .W22(W22TO24), .W23(W23TO24), .W24(W24TO24), .W25(W25TO24), .W26(W26TO24), .W27(W27TO24), .W28(W28TO24), .W29(W29TO24), .W30(W30TO24), .W31(W31TO24), .W32(W32TO24), .W33(W33TO24), .W34(W34TO24), .W35(W35TO24), .W36(W36TO24), .W37(W37TO24), .W38(W38TO24), .W39(W39TO24), .W40(W40TO24), .W41(W41TO24), .W42(W42TO24), .W43(W43TO24), .W44(W44TO24), .W45(W45TO24), .W46(W46TO24), .W47(W47TO24), .W48(W48TO24), .W49(W49TO24), .W50(W50TO24), .W51(W51TO24), .W52(W52TO24), .W53(W53TO24), .W54(W54TO24), .W55(W55TO24), .W56(W56TO24), .W57(W57TO24), .W58(W58TO24), .W59(W59TO24), .W60(W60TO24), .W61(W61TO24), .W62(W62TO24), .W63(W63TO24), .W64(W64TO24)) neuron24(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out24));
neuron65in #(.BIAS(BIAS25), .W0(W0TO25), .W1(W1TO25), .W2(W2TO25), .W3(W3TO25), .W4(W4TO25), .W5(W5TO25), .W6(W6TO25), .W7(W7TO25), .W8(W8TO25), .W9(W9TO25), .W10(W10TO25), .W11(W11TO25), .W12(W12TO25), .W13(W13TO25), .W14(W14TO25), .W15(W15TO25), .W16(W16TO25), .W17(W17TO25), .W18(W18TO25), .W19(W19TO25), .W20(W20TO25), .W21(W21TO25), .W22(W22TO25), .W23(W23TO25), .W24(W24TO25), .W25(W25TO25), .W26(W26TO25), .W27(W27TO25), .W28(W28TO25), .W29(W29TO25), .W30(W30TO25), .W31(W31TO25), .W32(W32TO25), .W33(W33TO25), .W34(W34TO25), .W35(W35TO25), .W36(W36TO25), .W37(W37TO25), .W38(W38TO25), .W39(W39TO25), .W40(W40TO25), .W41(W41TO25), .W42(W42TO25), .W43(W43TO25), .W44(W44TO25), .W45(W45TO25), .W46(W46TO25), .W47(W47TO25), .W48(W48TO25), .W49(W49TO25), .W50(W50TO25), .W51(W51TO25), .W52(W52TO25), .W53(W53TO25), .W54(W54TO25), .W55(W55TO25), .W56(W56TO25), .W57(W57TO25), .W58(W58TO25), .W59(W59TO25), .W60(W60TO25), .W61(W61TO25), .W62(W62TO25), .W63(W63TO25), .W64(W64TO25)) neuron25(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out25));
neuron65in #(.BIAS(BIAS26), .W0(W0TO26), .W1(W1TO26), .W2(W2TO26), .W3(W3TO26), .W4(W4TO26), .W5(W5TO26), .W6(W6TO26), .W7(W7TO26), .W8(W8TO26), .W9(W9TO26), .W10(W10TO26), .W11(W11TO26), .W12(W12TO26), .W13(W13TO26), .W14(W14TO26), .W15(W15TO26), .W16(W16TO26), .W17(W17TO26), .W18(W18TO26), .W19(W19TO26), .W20(W20TO26), .W21(W21TO26), .W22(W22TO26), .W23(W23TO26), .W24(W24TO26), .W25(W25TO26), .W26(W26TO26), .W27(W27TO26), .W28(W28TO26), .W29(W29TO26), .W30(W30TO26), .W31(W31TO26), .W32(W32TO26), .W33(W33TO26), .W34(W34TO26), .W35(W35TO26), .W36(W36TO26), .W37(W37TO26), .W38(W38TO26), .W39(W39TO26), .W40(W40TO26), .W41(W41TO26), .W42(W42TO26), .W43(W43TO26), .W44(W44TO26), .W45(W45TO26), .W46(W46TO26), .W47(W47TO26), .W48(W48TO26), .W49(W49TO26), .W50(W50TO26), .W51(W51TO26), .W52(W52TO26), .W53(W53TO26), .W54(W54TO26), .W55(W55TO26), .W56(W56TO26), .W57(W57TO26), .W58(W58TO26), .W59(W59TO26), .W60(W60TO26), .W61(W61TO26), .W62(W62TO26), .W63(W63TO26), .W64(W64TO26)) neuron26(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out26));
neuron65in #(.BIAS(BIAS27), .W0(W0TO27), .W1(W1TO27), .W2(W2TO27), .W3(W3TO27), .W4(W4TO27), .W5(W5TO27), .W6(W6TO27), .W7(W7TO27), .W8(W8TO27), .W9(W9TO27), .W10(W10TO27), .W11(W11TO27), .W12(W12TO27), .W13(W13TO27), .W14(W14TO27), .W15(W15TO27), .W16(W16TO27), .W17(W17TO27), .W18(W18TO27), .W19(W19TO27), .W20(W20TO27), .W21(W21TO27), .W22(W22TO27), .W23(W23TO27), .W24(W24TO27), .W25(W25TO27), .W26(W26TO27), .W27(W27TO27), .W28(W28TO27), .W29(W29TO27), .W30(W30TO27), .W31(W31TO27), .W32(W32TO27), .W33(W33TO27), .W34(W34TO27), .W35(W35TO27), .W36(W36TO27), .W37(W37TO27), .W38(W38TO27), .W39(W39TO27), .W40(W40TO27), .W41(W41TO27), .W42(W42TO27), .W43(W43TO27), .W44(W44TO27), .W45(W45TO27), .W46(W46TO27), .W47(W47TO27), .W48(W48TO27), .W49(W49TO27), .W50(W50TO27), .W51(W51TO27), .W52(W52TO27), .W53(W53TO27), .W54(W54TO27), .W55(W55TO27), .W56(W56TO27), .W57(W57TO27), .W58(W58TO27), .W59(W59TO27), .W60(W60TO27), .W61(W61TO27), .W62(W62TO27), .W63(W63TO27), .W64(W64TO27)) neuron27(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out27));
neuron65in #(.BIAS(BIAS28), .W0(W0TO28), .W1(W1TO28), .W2(W2TO28), .W3(W3TO28), .W4(W4TO28), .W5(W5TO28), .W6(W6TO28), .W7(W7TO28), .W8(W8TO28), .W9(W9TO28), .W10(W10TO28), .W11(W11TO28), .W12(W12TO28), .W13(W13TO28), .W14(W14TO28), .W15(W15TO28), .W16(W16TO28), .W17(W17TO28), .W18(W18TO28), .W19(W19TO28), .W20(W20TO28), .W21(W21TO28), .W22(W22TO28), .W23(W23TO28), .W24(W24TO28), .W25(W25TO28), .W26(W26TO28), .W27(W27TO28), .W28(W28TO28), .W29(W29TO28), .W30(W30TO28), .W31(W31TO28), .W32(W32TO28), .W33(W33TO28), .W34(W34TO28), .W35(W35TO28), .W36(W36TO28), .W37(W37TO28), .W38(W38TO28), .W39(W39TO28), .W40(W40TO28), .W41(W41TO28), .W42(W42TO28), .W43(W43TO28), .W44(W44TO28), .W45(W45TO28), .W46(W46TO28), .W47(W47TO28), .W48(W48TO28), .W49(W49TO28), .W50(W50TO28), .W51(W51TO28), .W52(W52TO28), .W53(W53TO28), .W54(W54TO28), .W55(W55TO28), .W56(W56TO28), .W57(W57TO28), .W58(W58TO28), .W59(W59TO28), .W60(W60TO28), .W61(W61TO28), .W62(W62TO28), .W63(W63TO28), .W64(W64TO28)) neuron28(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out28));
neuron65in #(.BIAS(BIAS29), .W0(W0TO29), .W1(W1TO29), .W2(W2TO29), .W3(W3TO29), .W4(W4TO29), .W5(W5TO29), .W6(W6TO29), .W7(W7TO29), .W8(W8TO29), .W9(W9TO29), .W10(W10TO29), .W11(W11TO29), .W12(W12TO29), .W13(W13TO29), .W14(W14TO29), .W15(W15TO29), .W16(W16TO29), .W17(W17TO29), .W18(W18TO29), .W19(W19TO29), .W20(W20TO29), .W21(W21TO29), .W22(W22TO29), .W23(W23TO29), .W24(W24TO29), .W25(W25TO29), .W26(W26TO29), .W27(W27TO29), .W28(W28TO29), .W29(W29TO29), .W30(W30TO29), .W31(W31TO29), .W32(W32TO29), .W33(W33TO29), .W34(W34TO29), .W35(W35TO29), .W36(W36TO29), .W37(W37TO29), .W38(W38TO29), .W39(W39TO29), .W40(W40TO29), .W41(W41TO29), .W42(W42TO29), .W43(W43TO29), .W44(W44TO29), .W45(W45TO29), .W46(W46TO29), .W47(W47TO29), .W48(W48TO29), .W49(W49TO29), .W50(W50TO29), .W51(W51TO29), .W52(W52TO29), .W53(W53TO29), .W54(W54TO29), .W55(W55TO29), .W56(W56TO29), .W57(W57TO29), .W58(W58TO29), .W59(W59TO29), .W60(W60TO29), .W61(W61TO29), .W62(W62TO29), .W63(W63TO29), .W64(W64TO29)) neuron29(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out29));
neuron65in #(.BIAS(BIAS30), .W0(W0TO30), .W1(W1TO30), .W2(W2TO30), .W3(W3TO30), .W4(W4TO30), .W5(W5TO30), .W6(W6TO30), .W7(W7TO30), .W8(W8TO30), .W9(W9TO30), .W10(W10TO30), .W11(W11TO30), .W12(W12TO30), .W13(W13TO30), .W14(W14TO30), .W15(W15TO30), .W16(W16TO30), .W17(W17TO30), .W18(W18TO30), .W19(W19TO30), .W20(W20TO30), .W21(W21TO30), .W22(W22TO30), .W23(W23TO30), .W24(W24TO30), .W25(W25TO30), .W26(W26TO30), .W27(W27TO30), .W28(W28TO30), .W29(W29TO30), .W30(W30TO30), .W31(W31TO30), .W32(W32TO30), .W33(W33TO30), .W34(W34TO30), .W35(W35TO30), .W36(W36TO30), .W37(W37TO30), .W38(W38TO30), .W39(W39TO30), .W40(W40TO30), .W41(W41TO30), .W42(W42TO30), .W43(W43TO30), .W44(W44TO30), .W45(W45TO30), .W46(W46TO30), .W47(W47TO30), .W48(W48TO30), .W49(W49TO30), .W50(W50TO30), .W51(W51TO30), .W52(W52TO30), .W53(W53TO30), .W54(W54TO30), .W55(W55TO30), .W56(W56TO30), .W57(W57TO30), .W58(W58TO30), .W59(W59TO30), .W60(W60TO30), .W61(W61TO30), .W62(W62TO30), .W63(W63TO30), .W64(W64TO30)) neuron30(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out30));
neuron65in #(.BIAS(BIAS31), .W0(W0TO31), .W1(W1TO31), .W2(W2TO31), .W3(W3TO31), .W4(W4TO31), .W5(W5TO31), .W6(W6TO31), .W7(W7TO31), .W8(W8TO31), .W9(W9TO31), .W10(W10TO31), .W11(W11TO31), .W12(W12TO31), .W13(W13TO31), .W14(W14TO31), .W15(W15TO31), .W16(W16TO31), .W17(W17TO31), .W18(W18TO31), .W19(W19TO31), .W20(W20TO31), .W21(W21TO31), .W22(W22TO31), .W23(W23TO31), .W24(W24TO31), .W25(W25TO31), .W26(W26TO31), .W27(W27TO31), .W28(W28TO31), .W29(W29TO31), .W30(W30TO31), .W31(W31TO31), .W32(W32TO31), .W33(W33TO31), .W34(W34TO31), .W35(W35TO31), .W36(W36TO31), .W37(W37TO31), .W38(W38TO31), .W39(W39TO31), .W40(W40TO31), .W41(W41TO31), .W42(W42TO31), .W43(W43TO31), .W44(W44TO31), .W45(W45TO31), .W46(W46TO31), .W47(W47TO31), .W48(W48TO31), .W49(W49TO31), .W50(W50TO31), .W51(W51TO31), .W52(W52TO31), .W53(W53TO31), .W54(W54TO31), .W55(W55TO31), .W56(W56TO31), .W57(W57TO31), .W58(W58TO31), .W59(W59TO31), .W60(W60TO31), .W61(W61TO31), .W62(W62TO31), .W63(W63TO31), .W64(W64TO31)) neuron31(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out31));
neuron65in #(.BIAS(BIAS32), .W0(W0TO32), .W1(W1TO32), .W2(W2TO32), .W3(W3TO32), .W4(W4TO32), .W5(W5TO32), .W6(W6TO32), .W7(W7TO32), .W8(W8TO32), .W9(W9TO32), .W10(W10TO32), .W11(W11TO32), .W12(W12TO32), .W13(W13TO32), .W14(W14TO32), .W15(W15TO32), .W16(W16TO32), .W17(W17TO32), .W18(W18TO32), .W19(W19TO32), .W20(W20TO32), .W21(W21TO32), .W22(W22TO32), .W23(W23TO32), .W24(W24TO32), .W25(W25TO32), .W26(W26TO32), .W27(W27TO32), .W28(W28TO32), .W29(W29TO32), .W30(W30TO32), .W31(W31TO32), .W32(W32TO32), .W33(W33TO32), .W34(W34TO32), .W35(W35TO32), .W36(W36TO32), .W37(W37TO32), .W38(W38TO32), .W39(W39TO32), .W40(W40TO32), .W41(W41TO32), .W42(W42TO32), .W43(W43TO32), .W44(W44TO32), .W45(W45TO32), .W46(W46TO32), .W47(W47TO32), .W48(W48TO32), .W49(W49TO32), .W50(W50TO32), .W51(W51TO32), .W52(W52TO32), .W53(W53TO32), .W54(W54TO32), .W55(W55TO32), .W56(W56TO32), .W57(W57TO32), .W58(W58TO32), .W59(W59TO32), .W60(W60TO32), .W61(W61TO32), .W62(W62TO32), .W63(W63TO32), .W64(W64TO32)) neuron32(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out32));
neuron65in #(.BIAS(BIAS33), .W0(W0TO33), .W1(W1TO33), .W2(W2TO33), .W3(W3TO33), .W4(W4TO33), .W5(W5TO33), .W6(W6TO33), .W7(W7TO33), .W8(W8TO33), .W9(W9TO33), .W10(W10TO33), .W11(W11TO33), .W12(W12TO33), .W13(W13TO33), .W14(W14TO33), .W15(W15TO33), .W16(W16TO33), .W17(W17TO33), .W18(W18TO33), .W19(W19TO33), .W20(W20TO33), .W21(W21TO33), .W22(W22TO33), .W23(W23TO33), .W24(W24TO33), .W25(W25TO33), .W26(W26TO33), .W27(W27TO33), .W28(W28TO33), .W29(W29TO33), .W30(W30TO33), .W31(W31TO33), .W32(W32TO33), .W33(W33TO33), .W34(W34TO33), .W35(W35TO33), .W36(W36TO33), .W37(W37TO33), .W38(W38TO33), .W39(W39TO33), .W40(W40TO33), .W41(W41TO33), .W42(W42TO33), .W43(W43TO33), .W44(W44TO33), .W45(W45TO33), .W46(W46TO33), .W47(W47TO33), .W48(W48TO33), .W49(W49TO33), .W50(W50TO33), .W51(W51TO33), .W52(W52TO33), .W53(W53TO33), .W54(W54TO33), .W55(W55TO33), .W56(W56TO33), .W57(W57TO33), .W58(W58TO33), .W59(W59TO33), .W60(W60TO33), .W61(W61TO33), .W62(W62TO33), .W63(W63TO33), .W64(W64TO33)) neuron33(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out33));
neuron65in #(.BIAS(BIAS34), .W0(W0TO34), .W1(W1TO34), .W2(W2TO34), .W3(W3TO34), .W4(W4TO34), .W5(W5TO34), .W6(W6TO34), .W7(W7TO34), .W8(W8TO34), .W9(W9TO34), .W10(W10TO34), .W11(W11TO34), .W12(W12TO34), .W13(W13TO34), .W14(W14TO34), .W15(W15TO34), .W16(W16TO34), .W17(W17TO34), .W18(W18TO34), .W19(W19TO34), .W20(W20TO34), .W21(W21TO34), .W22(W22TO34), .W23(W23TO34), .W24(W24TO34), .W25(W25TO34), .W26(W26TO34), .W27(W27TO34), .W28(W28TO34), .W29(W29TO34), .W30(W30TO34), .W31(W31TO34), .W32(W32TO34), .W33(W33TO34), .W34(W34TO34), .W35(W35TO34), .W36(W36TO34), .W37(W37TO34), .W38(W38TO34), .W39(W39TO34), .W40(W40TO34), .W41(W41TO34), .W42(W42TO34), .W43(W43TO34), .W44(W44TO34), .W45(W45TO34), .W46(W46TO34), .W47(W47TO34), .W48(W48TO34), .W49(W49TO34), .W50(W50TO34), .W51(W51TO34), .W52(W52TO34), .W53(W53TO34), .W54(W54TO34), .W55(W55TO34), .W56(W56TO34), .W57(W57TO34), .W58(W58TO34), .W59(W59TO34), .W60(W60TO34), .W61(W61TO34), .W62(W62TO34), .W63(W63TO34), .W64(W64TO34)) neuron34(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out34));
neuron65in #(.BIAS(BIAS35), .W0(W0TO35), .W1(W1TO35), .W2(W2TO35), .W3(W3TO35), .W4(W4TO35), .W5(W5TO35), .W6(W6TO35), .W7(W7TO35), .W8(W8TO35), .W9(W9TO35), .W10(W10TO35), .W11(W11TO35), .W12(W12TO35), .W13(W13TO35), .W14(W14TO35), .W15(W15TO35), .W16(W16TO35), .W17(W17TO35), .W18(W18TO35), .W19(W19TO35), .W20(W20TO35), .W21(W21TO35), .W22(W22TO35), .W23(W23TO35), .W24(W24TO35), .W25(W25TO35), .W26(W26TO35), .W27(W27TO35), .W28(W28TO35), .W29(W29TO35), .W30(W30TO35), .W31(W31TO35), .W32(W32TO35), .W33(W33TO35), .W34(W34TO35), .W35(W35TO35), .W36(W36TO35), .W37(W37TO35), .W38(W38TO35), .W39(W39TO35), .W40(W40TO35), .W41(W41TO35), .W42(W42TO35), .W43(W43TO35), .W44(W44TO35), .W45(W45TO35), .W46(W46TO35), .W47(W47TO35), .W48(W48TO35), .W49(W49TO35), .W50(W50TO35), .W51(W51TO35), .W52(W52TO35), .W53(W53TO35), .W54(W54TO35), .W55(W55TO35), .W56(W56TO35), .W57(W57TO35), .W58(W58TO35), .W59(W59TO35), .W60(W60TO35), .W61(W61TO35), .W62(W62TO35), .W63(W63TO35), .W64(W64TO35)) neuron35(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out35));
neuron65in #(.BIAS(BIAS36), .W0(W0TO36), .W1(W1TO36), .W2(W2TO36), .W3(W3TO36), .W4(W4TO36), .W5(W5TO36), .W6(W6TO36), .W7(W7TO36), .W8(W8TO36), .W9(W9TO36), .W10(W10TO36), .W11(W11TO36), .W12(W12TO36), .W13(W13TO36), .W14(W14TO36), .W15(W15TO36), .W16(W16TO36), .W17(W17TO36), .W18(W18TO36), .W19(W19TO36), .W20(W20TO36), .W21(W21TO36), .W22(W22TO36), .W23(W23TO36), .W24(W24TO36), .W25(W25TO36), .W26(W26TO36), .W27(W27TO36), .W28(W28TO36), .W29(W29TO36), .W30(W30TO36), .W31(W31TO36), .W32(W32TO36), .W33(W33TO36), .W34(W34TO36), .W35(W35TO36), .W36(W36TO36), .W37(W37TO36), .W38(W38TO36), .W39(W39TO36), .W40(W40TO36), .W41(W41TO36), .W42(W42TO36), .W43(W43TO36), .W44(W44TO36), .W45(W45TO36), .W46(W46TO36), .W47(W47TO36), .W48(W48TO36), .W49(W49TO36), .W50(W50TO36), .W51(W51TO36), .W52(W52TO36), .W53(W53TO36), .W54(W54TO36), .W55(W55TO36), .W56(W56TO36), .W57(W57TO36), .W58(W58TO36), .W59(W59TO36), .W60(W60TO36), .W61(W61TO36), .W62(W62TO36), .W63(W63TO36), .W64(W64TO36)) neuron36(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out36));
neuron65in #(.BIAS(BIAS37), .W0(W0TO37), .W1(W1TO37), .W2(W2TO37), .W3(W3TO37), .W4(W4TO37), .W5(W5TO37), .W6(W6TO37), .W7(W7TO37), .W8(W8TO37), .W9(W9TO37), .W10(W10TO37), .W11(W11TO37), .W12(W12TO37), .W13(W13TO37), .W14(W14TO37), .W15(W15TO37), .W16(W16TO37), .W17(W17TO37), .W18(W18TO37), .W19(W19TO37), .W20(W20TO37), .W21(W21TO37), .W22(W22TO37), .W23(W23TO37), .W24(W24TO37), .W25(W25TO37), .W26(W26TO37), .W27(W27TO37), .W28(W28TO37), .W29(W29TO37), .W30(W30TO37), .W31(W31TO37), .W32(W32TO37), .W33(W33TO37), .W34(W34TO37), .W35(W35TO37), .W36(W36TO37), .W37(W37TO37), .W38(W38TO37), .W39(W39TO37), .W40(W40TO37), .W41(W41TO37), .W42(W42TO37), .W43(W43TO37), .W44(W44TO37), .W45(W45TO37), .W46(W46TO37), .W47(W47TO37), .W48(W48TO37), .W49(W49TO37), .W50(W50TO37), .W51(W51TO37), .W52(W52TO37), .W53(W53TO37), .W54(W54TO37), .W55(W55TO37), .W56(W56TO37), .W57(W57TO37), .W58(W58TO37), .W59(W59TO37), .W60(W60TO37), .W61(W61TO37), .W62(W62TO37), .W63(W63TO37), .W64(W64TO37)) neuron37(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out37));
neuron65in #(.BIAS(BIAS38), .W0(W0TO38), .W1(W1TO38), .W2(W2TO38), .W3(W3TO38), .W4(W4TO38), .W5(W5TO38), .W6(W6TO38), .W7(W7TO38), .W8(W8TO38), .W9(W9TO38), .W10(W10TO38), .W11(W11TO38), .W12(W12TO38), .W13(W13TO38), .W14(W14TO38), .W15(W15TO38), .W16(W16TO38), .W17(W17TO38), .W18(W18TO38), .W19(W19TO38), .W20(W20TO38), .W21(W21TO38), .W22(W22TO38), .W23(W23TO38), .W24(W24TO38), .W25(W25TO38), .W26(W26TO38), .W27(W27TO38), .W28(W28TO38), .W29(W29TO38), .W30(W30TO38), .W31(W31TO38), .W32(W32TO38), .W33(W33TO38), .W34(W34TO38), .W35(W35TO38), .W36(W36TO38), .W37(W37TO38), .W38(W38TO38), .W39(W39TO38), .W40(W40TO38), .W41(W41TO38), .W42(W42TO38), .W43(W43TO38), .W44(W44TO38), .W45(W45TO38), .W46(W46TO38), .W47(W47TO38), .W48(W48TO38), .W49(W49TO38), .W50(W50TO38), .W51(W51TO38), .W52(W52TO38), .W53(W53TO38), .W54(W54TO38), .W55(W55TO38), .W56(W56TO38), .W57(W57TO38), .W58(W58TO38), .W59(W59TO38), .W60(W60TO38), .W61(W61TO38), .W62(W62TO38), .W63(W63TO38), .W64(W64TO38)) neuron38(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out38));
neuron65in #(.BIAS(BIAS39), .W0(W0TO39), .W1(W1TO39), .W2(W2TO39), .W3(W3TO39), .W4(W4TO39), .W5(W5TO39), .W6(W6TO39), .W7(W7TO39), .W8(W8TO39), .W9(W9TO39), .W10(W10TO39), .W11(W11TO39), .W12(W12TO39), .W13(W13TO39), .W14(W14TO39), .W15(W15TO39), .W16(W16TO39), .W17(W17TO39), .W18(W18TO39), .W19(W19TO39), .W20(W20TO39), .W21(W21TO39), .W22(W22TO39), .W23(W23TO39), .W24(W24TO39), .W25(W25TO39), .W26(W26TO39), .W27(W27TO39), .W28(W28TO39), .W29(W29TO39), .W30(W30TO39), .W31(W31TO39), .W32(W32TO39), .W33(W33TO39), .W34(W34TO39), .W35(W35TO39), .W36(W36TO39), .W37(W37TO39), .W38(W38TO39), .W39(W39TO39), .W40(W40TO39), .W41(W41TO39), .W42(W42TO39), .W43(W43TO39), .W44(W44TO39), .W45(W45TO39), .W46(W46TO39), .W47(W47TO39), .W48(W48TO39), .W49(W49TO39), .W50(W50TO39), .W51(W51TO39), .W52(W52TO39), .W53(W53TO39), .W54(W54TO39), .W55(W55TO39), .W56(W56TO39), .W57(W57TO39), .W58(W58TO39), .W59(W59TO39), .W60(W60TO39), .W61(W61TO39), .W62(W62TO39), .W63(W63TO39), .W64(W64TO39)) neuron39(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out39));
neuron65in #(.BIAS(BIAS40), .W0(W0TO40), .W1(W1TO40), .W2(W2TO40), .W3(W3TO40), .W4(W4TO40), .W5(W5TO40), .W6(W6TO40), .W7(W7TO40), .W8(W8TO40), .W9(W9TO40), .W10(W10TO40), .W11(W11TO40), .W12(W12TO40), .W13(W13TO40), .W14(W14TO40), .W15(W15TO40), .W16(W16TO40), .W17(W17TO40), .W18(W18TO40), .W19(W19TO40), .W20(W20TO40), .W21(W21TO40), .W22(W22TO40), .W23(W23TO40), .W24(W24TO40), .W25(W25TO40), .W26(W26TO40), .W27(W27TO40), .W28(W28TO40), .W29(W29TO40), .W30(W30TO40), .W31(W31TO40), .W32(W32TO40), .W33(W33TO40), .W34(W34TO40), .W35(W35TO40), .W36(W36TO40), .W37(W37TO40), .W38(W38TO40), .W39(W39TO40), .W40(W40TO40), .W41(W41TO40), .W42(W42TO40), .W43(W43TO40), .W44(W44TO40), .W45(W45TO40), .W46(W46TO40), .W47(W47TO40), .W48(W48TO40), .W49(W49TO40), .W50(W50TO40), .W51(W51TO40), .W52(W52TO40), .W53(W53TO40), .W54(W54TO40), .W55(W55TO40), .W56(W56TO40), .W57(W57TO40), .W58(W58TO40), .W59(W59TO40), .W60(W60TO40), .W61(W61TO40), .W62(W62TO40), .W63(W63TO40), .W64(W64TO40)) neuron40(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out40));
neuron65in #(.BIAS(BIAS41), .W0(W0TO41), .W1(W1TO41), .W2(W2TO41), .W3(W3TO41), .W4(W4TO41), .W5(W5TO41), .W6(W6TO41), .W7(W7TO41), .W8(W8TO41), .W9(W9TO41), .W10(W10TO41), .W11(W11TO41), .W12(W12TO41), .W13(W13TO41), .W14(W14TO41), .W15(W15TO41), .W16(W16TO41), .W17(W17TO41), .W18(W18TO41), .W19(W19TO41), .W20(W20TO41), .W21(W21TO41), .W22(W22TO41), .W23(W23TO41), .W24(W24TO41), .W25(W25TO41), .W26(W26TO41), .W27(W27TO41), .W28(W28TO41), .W29(W29TO41), .W30(W30TO41), .W31(W31TO41), .W32(W32TO41), .W33(W33TO41), .W34(W34TO41), .W35(W35TO41), .W36(W36TO41), .W37(W37TO41), .W38(W38TO41), .W39(W39TO41), .W40(W40TO41), .W41(W41TO41), .W42(W42TO41), .W43(W43TO41), .W44(W44TO41), .W45(W45TO41), .W46(W46TO41), .W47(W47TO41), .W48(W48TO41), .W49(W49TO41), .W50(W50TO41), .W51(W51TO41), .W52(W52TO41), .W53(W53TO41), .W54(W54TO41), .W55(W55TO41), .W56(W56TO41), .W57(W57TO41), .W58(W58TO41), .W59(W59TO41), .W60(W60TO41), .W61(W61TO41), .W62(W62TO41), .W63(W63TO41), .W64(W64TO41)) neuron41(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out41));
neuron65in #(.BIAS(BIAS42), .W0(W0TO42), .W1(W1TO42), .W2(W2TO42), .W3(W3TO42), .W4(W4TO42), .W5(W5TO42), .W6(W6TO42), .W7(W7TO42), .W8(W8TO42), .W9(W9TO42), .W10(W10TO42), .W11(W11TO42), .W12(W12TO42), .W13(W13TO42), .W14(W14TO42), .W15(W15TO42), .W16(W16TO42), .W17(W17TO42), .W18(W18TO42), .W19(W19TO42), .W20(W20TO42), .W21(W21TO42), .W22(W22TO42), .W23(W23TO42), .W24(W24TO42), .W25(W25TO42), .W26(W26TO42), .W27(W27TO42), .W28(W28TO42), .W29(W29TO42), .W30(W30TO42), .W31(W31TO42), .W32(W32TO42), .W33(W33TO42), .W34(W34TO42), .W35(W35TO42), .W36(W36TO42), .W37(W37TO42), .W38(W38TO42), .W39(W39TO42), .W40(W40TO42), .W41(W41TO42), .W42(W42TO42), .W43(W43TO42), .W44(W44TO42), .W45(W45TO42), .W46(W46TO42), .W47(W47TO42), .W48(W48TO42), .W49(W49TO42), .W50(W50TO42), .W51(W51TO42), .W52(W52TO42), .W53(W53TO42), .W54(W54TO42), .W55(W55TO42), .W56(W56TO42), .W57(W57TO42), .W58(W58TO42), .W59(W59TO42), .W60(W60TO42), .W61(W61TO42), .W62(W62TO42), .W63(W63TO42), .W64(W64TO42)) neuron42(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out42));
neuron65in #(.BIAS(BIAS43), .W0(W0TO43), .W1(W1TO43), .W2(W2TO43), .W3(W3TO43), .W4(W4TO43), .W5(W5TO43), .W6(W6TO43), .W7(W7TO43), .W8(W8TO43), .W9(W9TO43), .W10(W10TO43), .W11(W11TO43), .W12(W12TO43), .W13(W13TO43), .W14(W14TO43), .W15(W15TO43), .W16(W16TO43), .W17(W17TO43), .W18(W18TO43), .W19(W19TO43), .W20(W20TO43), .W21(W21TO43), .W22(W22TO43), .W23(W23TO43), .W24(W24TO43), .W25(W25TO43), .W26(W26TO43), .W27(W27TO43), .W28(W28TO43), .W29(W29TO43), .W30(W30TO43), .W31(W31TO43), .W32(W32TO43), .W33(W33TO43), .W34(W34TO43), .W35(W35TO43), .W36(W36TO43), .W37(W37TO43), .W38(W38TO43), .W39(W39TO43), .W40(W40TO43), .W41(W41TO43), .W42(W42TO43), .W43(W43TO43), .W44(W44TO43), .W45(W45TO43), .W46(W46TO43), .W47(W47TO43), .W48(W48TO43), .W49(W49TO43), .W50(W50TO43), .W51(W51TO43), .W52(W52TO43), .W53(W53TO43), .W54(W54TO43), .W55(W55TO43), .W56(W56TO43), .W57(W57TO43), .W58(W58TO43), .W59(W59TO43), .W60(W60TO43), .W61(W61TO43), .W62(W62TO43), .W63(W63TO43), .W64(W64TO43)) neuron43(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out43));
neuron65in #(.BIAS(BIAS44), .W0(W0TO44), .W1(W1TO44), .W2(W2TO44), .W3(W3TO44), .W4(W4TO44), .W5(W5TO44), .W6(W6TO44), .W7(W7TO44), .W8(W8TO44), .W9(W9TO44), .W10(W10TO44), .W11(W11TO44), .W12(W12TO44), .W13(W13TO44), .W14(W14TO44), .W15(W15TO44), .W16(W16TO44), .W17(W17TO44), .W18(W18TO44), .W19(W19TO44), .W20(W20TO44), .W21(W21TO44), .W22(W22TO44), .W23(W23TO44), .W24(W24TO44), .W25(W25TO44), .W26(W26TO44), .W27(W27TO44), .W28(W28TO44), .W29(W29TO44), .W30(W30TO44), .W31(W31TO44), .W32(W32TO44), .W33(W33TO44), .W34(W34TO44), .W35(W35TO44), .W36(W36TO44), .W37(W37TO44), .W38(W38TO44), .W39(W39TO44), .W40(W40TO44), .W41(W41TO44), .W42(W42TO44), .W43(W43TO44), .W44(W44TO44), .W45(W45TO44), .W46(W46TO44), .W47(W47TO44), .W48(W48TO44), .W49(W49TO44), .W50(W50TO44), .W51(W51TO44), .W52(W52TO44), .W53(W53TO44), .W54(W54TO44), .W55(W55TO44), .W56(W56TO44), .W57(W57TO44), .W58(W58TO44), .W59(W59TO44), .W60(W60TO44), .W61(W61TO44), .W62(W62TO44), .W63(W63TO44), .W64(W64TO44)) neuron44(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out44));
neuron65in #(.BIAS(BIAS45), .W0(W0TO45), .W1(W1TO45), .W2(W2TO45), .W3(W3TO45), .W4(W4TO45), .W5(W5TO45), .W6(W6TO45), .W7(W7TO45), .W8(W8TO45), .W9(W9TO45), .W10(W10TO45), .W11(W11TO45), .W12(W12TO45), .W13(W13TO45), .W14(W14TO45), .W15(W15TO45), .W16(W16TO45), .W17(W17TO45), .W18(W18TO45), .W19(W19TO45), .W20(W20TO45), .W21(W21TO45), .W22(W22TO45), .W23(W23TO45), .W24(W24TO45), .W25(W25TO45), .W26(W26TO45), .W27(W27TO45), .W28(W28TO45), .W29(W29TO45), .W30(W30TO45), .W31(W31TO45), .W32(W32TO45), .W33(W33TO45), .W34(W34TO45), .W35(W35TO45), .W36(W36TO45), .W37(W37TO45), .W38(W38TO45), .W39(W39TO45), .W40(W40TO45), .W41(W41TO45), .W42(W42TO45), .W43(W43TO45), .W44(W44TO45), .W45(W45TO45), .W46(W46TO45), .W47(W47TO45), .W48(W48TO45), .W49(W49TO45), .W50(W50TO45), .W51(W51TO45), .W52(W52TO45), .W53(W53TO45), .W54(W54TO45), .W55(W55TO45), .W56(W56TO45), .W57(W57TO45), .W58(W58TO45), .W59(W59TO45), .W60(W60TO45), .W61(W61TO45), .W62(W62TO45), .W63(W63TO45), .W64(W64TO45)) neuron45(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out45));
neuron65in #(.BIAS(BIAS46), .W0(W0TO46), .W1(W1TO46), .W2(W2TO46), .W3(W3TO46), .W4(W4TO46), .W5(W5TO46), .W6(W6TO46), .W7(W7TO46), .W8(W8TO46), .W9(W9TO46), .W10(W10TO46), .W11(W11TO46), .W12(W12TO46), .W13(W13TO46), .W14(W14TO46), .W15(W15TO46), .W16(W16TO46), .W17(W17TO46), .W18(W18TO46), .W19(W19TO46), .W20(W20TO46), .W21(W21TO46), .W22(W22TO46), .W23(W23TO46), .W24(W24TO46), .W25(W25TO46), .W26(W26TO46), .W27(W27TO46), .W28(W28TO46), .W29(W29TO46), .W30(W30TO46), .W31(W31TO46), .W32(W32TO46), .W33(W33TO46), .W34(W34TO46), .W35(W35TO46), .W36(W36TO46), .W37(W37TO46), .W38(W38TO46), .W39(W39TO46), .W40(W40TO46), .W41(W41TO46), .W42(W42TO46), .W43(W43TO46), .W44(W44TO46), .W45(W45TO46), .W46(W46TO46), .W47(W47TO46), .W48(W48TO46), .W49(W49TO46), .W50(W50TO46), .W51(W51TO46), .W52(W52TO46), .W53(W53TO46), .W54(W54TO46), .W55(W55TO46), .W56(W56TO46), .W57(W57TO46), .W58(W58TO46), .W59(W59TO46), .W60(W60TO46), .W61(W61TO46), .W62(W62TO46), .W63(W63TO46), .W64(W64TO46)) neuron46(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out46));
neuron65in #(.BIAS(BIAS47), .W0(W0TO47), .W1(W1TO47), .W2(W2TO47), .W3(W3TO47), .W4(W4TO47), .W5(W5TO47), .W6(W6TO47), .W7(W7TO47), .W8(W8TO47), .W9(W9TO47), .W10(W10TO47), .W11(W11TO47), .W12(W12TO47), .W13(W13TO47), .W14(W14TO47), .W15(W15TO47), .W16(W16TO47), .W17(W17TO47), .W18(W18TO47), .W19(W19TO47), .W20(W20TO47), .W21(W21TO47), .W22(W22TO47), .W23(W23TO47), .W24(W24TO47), .W25(W25TO47), .W26(W26TO47), .W27(W27TO47), .W28(W28TO47), .W29(W29TO47), .W30(W30TO47), .W31(W31TO47), .W32(W32TO47), .W33(W33TO47), .W34(W34TO47), .W35(W35TO47), .W36(W36TO47), .W37(W37TO47), .W38(W38TO47), .W39(W39TO47), .W40(W40TO47), .W41(W41TO47), .W42(W42TO47), .W43(W43TO47), .W44(W44TO47), .W45(W45TO47), .W46(W46TO47), .W47(W47TO47), .W48(W48TO47), .W49(W49TO47), .W50(W50TO47), .W51(W51TO47), .W52(W52TO47), .W53(W53TO47), .W54(W54TO47), .W55(W55TO47), .W56(W56TO47), .W57(W57TO47), .W58(W58TO47), .W59(W59TO47), .W60(W60TO47), .W61(W61TO47), .W62(W62TO47), .W63(W63TO47), .W64(W64TO47)) neuron47(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out47));
neuron65in #(.BIAS(BIAS48), .W0(W0TO48), .W1(W1TO48), .W2(W2TO48), .W3(W3TO48), .W4(W4TO48), .W5(W5TO48), .W6(W6TO48), .W7(W7TO48), .W8(W8TO48), .W9(W9TO48), .W10(W10TO48), .W11(W11TO48), .W12(W12TO48), .W13(W13TO48), .W14(W14TO48), .W15(W15TO48), .W16(W16TO48), .W17(W17TO48), .W18(W18TO48), .W19(W19TO48), .W20(W20TO48), .W21(W21TO48), .W22(W22TO48), .W23(W23TO48), .W24(W24TO48), .W25(W25TO48), .W26(W26TO48), .W27(W27TO48), .W28(W28TO48), .W29(W29TO48), .W30(W30TO48), .W31(W31TO48), .W32(W32TO48), .W33(W33TO48), .W34(W34TO48), .W35(W35TO48), .W36(W36TO48), .W37(W37TO48), .W38(W38TO48), .W39(W39TO48), .W40(W40TO48), .W41(W41TO48), .W42(W42TO48), .W43(W43TO48), .W44(W44TO48), .W45(W45TO48), .W46(W46TO48), .W47(W47TO48), .W48(W48TO48), .W49(W49TO48), .W50(W50TO48), .W51(W51TO48), .W52(W52TO48), .W53(W53TO48), .W54(W54TO48), .W55(W55TO48), .W56(W56TO48), .W57(W57TO48), .W58(W58TO48), .W59(W59TO48), .W60(W60TO48), .W61(W61TO48), .W62(W62TO48), .W63(W63TO48), .W64(W64TO48)) neuron48(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out48));
neuron65in #(.BIAS(BIAS49), .W0(W0TO49), .W1(W1TO49), .W2(W2TO49), .W3(W3TO49), .W4(W4TO49), .W5(W5TO49), .W6(W6TO49), .W7(W7TO49), .W8(W8TO49), .W9(W9TO49), .W10(W10TO49), .W11(W11TO49), .W12(W12TO49), .W13(W13TO49), .W14(W14TO49), .W15(W15TO49), .W16(W16TO49), .W17(W17TO49), .W18(W18TO49), .W19(W19TO49), .W20(W20TO49), .W21(W21TO49), .W22(W22TO49), .W23(W23TO49), .W24(W24TO49), .W25(W25TO49), .W26(W26TO49), .W27(W27TO49), .W28(W28TO49), .W29(W29TO49), .W30(W30TO49), .W31(W31TO49), .W32(W32TO49), .W33(W33TO49), .W34(W34TO49), .W35(W35TO49), .W36(W36TO49), .W37(W37TO49), .W38(W38TO49), .W39(W39TO49), .W40(W40TO49), .W41(W41TO49), .W42(W42TO49), .W43(W43TO49), .W44(W44TO49), .W45(W45TO49), .W46(W46TO49), .W47(W47TO49), .W48(W48TO49), .W49(W49TO49), .W50(W50TO49), .W51(W51TO49), .W52(W52TO49), .W53(W53TO49), .W54(W54TO49), .W55(W55TO49), .W56(W56TO49), .W57(W57TO49), .W58(W58TO49), .W59(W59TO49), .W60(W60TO49), .W61(W61TO49), .W62(W62TO49), .W63(W63TO49), .W64(W64TO49)) neuron49(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out49));
neuron65in #(.BIAS(BIAS50), .W0(W0TO50), .W1(W1TO50), .W2(W2TO50), .W3(W3TO50), .W4(W4TO50), .W5(W5TO50), .W6(W6TO50), .W7(W7TO50), .W8(W8TO50), .W9(W9TO50), .W10(W10TO50), .W11(W11TO50), .W12(W12TO50), .W13(W13TO50), .W14(W14TO50), .W15(W15TO50), .W16(W16TO50), .W17(W17TO50), .W18(W18TO50), .W19(W19TO50), .W20(W20TO50), .W21(W21TO50), .W22(W22TO50), .W23(W23TO50), .W24(W24TO50), .W25(W25TO50), .W26(W26TO50), .W27(W27TO50), .W28(W28TO50), .W29(W29TO50), .W30(W30TO50), .W31(W31TO50), .W32(W32TO50), .W33(W33TO50), .W34(W34TO50), .W35(W35TO50), .W36(W36TO50), .W37(W37TO50), .W38(W38TO50), .W39(W39TO50), .W40(W40TO50), .W41(W41TO50), .W42(W42TO50), .W43(W43TO50), .W44(W44TO50), .W45(W45TO50), .W46(W46TO50), .W47(W47TO50), .W48(W48TO50), .W49(W49TO50), .W50(W50TO50), .W51(W51TO50), .W52(W52TO50), .W53(W53TO50), .W54(W54TO50), .W55(W55TO50), .W56(W56TO50), .W57(W57TO50), .W58(W58TO50), .W59(W59TO50), .W60(W60TO50), .W61(W61TO50), .W62(W62TO50), .W63(W63TO50), .W64(W64TO50)) neuron50(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out50));
neuron65in #(.BIAS(BIAS51), .W0(W0TO51), .W1(W1TO51), .W2(W2TO51), .W3(W3TO51), .W4(W4TO51), .W5(W5TO51), .W6(W6TO51), .W7(W7TO51), .W8(W8TO51), .W9(W9TO51), .W10(W10TO51), .W11(W11TO51), .W12(W12TO51), .W13(W13TO51), .W14(W14TO51), .W15(W15TO51), .W16(W16TO51), .W17(W17TO51), .W18(W18TO51), .W19(W19TO51), .W20(W20TO51), .W21(W21TO51), .W22(W22TO51), .W23(W23TO51), .W24(W24TO51), .W25(W25TO51), .W26(W26TO51), .W27(W27TO51), .W28(W28TO51), .W29(W29TO51), .W30(W30TO51), .W31(W31TO51), .W32(W32TO51), .W33(W33TO51), .W34(W34TO51), .W35(W35TO51), .W36(W36TO51), .W37(W37TO51), .W38(W38TO51), .W39(W39TO51), .W40(W40TO51), .W41(W41TO51), .W42(W42TO51), .W43(W43TO51), .W44(W44TO51), .W45(W45TO51), .W46(W46TO51), .W47(W47TO51), .W48(W48TO51), .W49(W49TO51), .W50(W50TO51), .W51(W51TO51), .W52(W52TO51), .W53(W53TO51), .W54(W54TO51), .W55(W55TO51), .W56(W56TO51), .W57(W57TO51), .W58(W58TO51), .W59(W59TO51), .W60(W60TO51), .W61(W61TO51), .W62(W62TO51), .W63(W63TO51), .W64(W64TO51)) neuron51(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out51));
neuron65in #(.BIAS(BIAS52), .W0(W0TO52), .W1(W1TO52), .W2(W2TO52), .W3(W3TO52), .W4(W4TO52), .W5(W5TO52), .W6(W6TO52), .W7(W7TO52), .W8(W8TO52), .W9(W9TO52), .W10(W10TO52), .W11(W11TO52), .W12(W12TO52), .W13(W13TO52), .W14(W14TO52), .W15(W15TO52), .W16(W16TO52), .W17(W17TO52), .W18(W18TO52), .W19(W19TO52), .W20(W20TO52), .W21(W21TO52), .W22(W22TO52), .W23(W23TO52), .W24(W24TO52), .W25(W25TO52), .W26(W26TO52), .W27(W27TO52), .W28(W28TO52), .W29(W29TO52), .W30(W30TO52), .W31(W31TO52), .W32(W32TO52), .W33(W33TO52), .W34(W34TO52), .W35(W35TO52), .W36(W36TO52), .W37(W37TO52), .W38(W38TO52), .W39(W39TO52), .W40(W40TO52), .W41(W41TO52), .W42(W42TO52), .W43(W43TO52), .W44(W44TO52), .W45(W45TO52), .W46(W46TO52), .W47(W47TO52), .W48(W48TO52), .W49(W49TO52), .W50(W50TO52), .W51(W51TO52), .W52(W52TO52), .W53(W53TO52), .W54(W54TO52), .W55(W55TO52), .W56(W56TO52), .W57(W57TO52), .W58(W58TO52), .W59(W59TO52), .W60(W60TO52), .W61(W61TO52), .W62(W62TO52), .W63(W63TO52), .W64(W64TO52)) neuron52(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out52));
neuron65in #(.BIAS(BIAS53), .W0(W0TO53), .W1(W1TO53), .W2(W2TO53), .W3(W3TO53), .W4(W4TO53), .W5(W5TO53), .W6(W6TO53), .W7(W7TO53), .W8(W8TO53), .W9(W9TO53), .W10(W10TO53), .W11(W11TO53), .W12(W12TO53), .W13(W13TO53), .W14(W14TO53), .W15(W15TO53), .W16(W16TO53), .W17(W17TO53), .W18(W18TO53), .W19(W19TO53), .W20(W20TO53), .W21(W21TO53), .W22(W22TO53), .W23(W23TO53), .W24(W24TO53), .W25(W25TO53), .W26(W26TO53), .W27(W27TO53), .W28(W28TO53), .W29(W29TO53), .W30(W30TO53), .W31(W31TO53), .W32(W32TO53), .W33(W33TO53), .W34(W34TO53), .W35(W35TO53), .W36(W36TO53), .W37(W37TO53), .W38(W38TO53), .W39(W39TO53), .W40(W40TO53), .W41(W41TO53), .W42(W42TO53), .W43(W43TO53), .W44(W44TO53), .W45(W45TO53), .W46(W46TO53), .W47(W47TO53), .W48(W48TO53), .W49(W49TO53), .W50(W50TO53), .W51(W51TO53), .W52(W52TO53), .W53(W53TO53), .W54(W54TO53), .W55(W55TO53), .W56(W56TO53), .W57(W57TO53), .W58(W58TO53), .W59(W59TO53), .W60(W60TO53), .W61(W61TO53), .W62(W62TO53), .W63(W63TO53), .W64(W64TO53)) neuron53(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out53));
neuron65in #(.BIAS(BIAS54), .W0(W0TO54), .W1(W1TO54), .W2(W2TO54), .W3(W3TO54), .W4(W4TO54), .W5(W5TO54), .W6(W6TO54), .W7(W7TO54), .W8(W8TO54), .W9(W9TO54), .W10(W10TO54), .W11(W11TO54), .W12(W12TO54), .W13(W13TO54), .W14(W14TO54), .W15(W15TO54), .W16(W16TO54), .W17(W17TO54), .W18(W18TO54), .W19(W19TO54), .W20(W20TO54), .W21(W21TO54), .W22(W22TO54), .W23(W23TO54), .W24(W24TO54), .W25(W25TO54), .W26(W26TO54), .W27(W27TO54), .W28(W28TO54), .W29(W29TO54), .W30(W30TO54), .W31(W31TO54), .W32(W32TO54), .W33(W33TO54), .W34(W34TO54), .W35(W35TO54), .W36(W36TO54), .W37(W37TO54), .W38(W38TO54), .W39(W39TO54), .W40(W40TO54), .W41(W41TO54), .W42(W42TO54), .W43(W43TO54), .W44(W44TO54), .W45(W45TO54), .W46(W46TO54), .W47(W47TO54), .W48(W48TO54), .W49(W49TO54), .W50(W50TO54), .W51(W51TO54), .W52(W52TO54), .W53(W53TO54), .W54(W54TO54), .W55(W55TO54), .W56(W56TO54), .W57(W57TO54), .W58(W58TO54), .W59(W59TO54), .W60(W60TO54), .W61(W61TO54), .W62(W62TO54), .W63(W63TO54), .W64(W64TO54)) neuron54(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out54));
neuron65in #(.BIAS(BIAS55), .W0(W0TO55), .W1(W1TO55), .W2(W2TO55), .W3(W3TO55), .W4(W4TO55), .W5(W5TO55), .W6(W6TO55), .W7(W7TO55), .W8(W8TO55), .W9(W9TO55), .W10(W10TO55), .W11(W11TO55), .W12(W12TO55), .W13(W13TO55), .W14(W14TO55), .W15(W15TO55), .W16(W16TO55), .W17(W17TO55), .W18(W18TO55), .W19(W19TO55), .W20(W20TO55), .W21(W21TO55), .W22(W22TO55), .W23(W23TO55), .W24(W24TO55), .W25(W25TO55), .W26(W26TO55), .W27(W27TO55), .W28(W28TO55), .W29(W29TO55), .W30(W30TO55), .W31(W31TO55), .W32(W32TO55), .W33(W33TO55), .W34(W34TO55), .W35(W35TO55), .W36(W36TO55), .W37(W37TO55), .W38(W38TO55), .W39(W39TO55), .W40(W40TO55), .W41(W41TO55), .W42(W42TO55), .W43(W43TO55), .W44(W44TO55), .W45(W45TO55), .W46(W46TO55), .W47(W47TO55), .W48(W48TO55), .W49(W49TO55), .W50(W50TO55), .W51(W51TO55), .W52(W52TO55), .W53(W53TO55), .W54(W54TO55), .W55(W55TO55), .W56(W56TO55), .W57(W57TO55), .W58(W58TO55), .W59(W59TO55), .W60(W60TO55), .W61(W61TO55), .W62(W62TO55), .W63(W63TO55), .W64(W64TO55)) neuron55(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out55));
neuron65in #(.BIAS(BIAS56), .W0(W0TO56), .W1(W1TO56), .W2(W2TO56), .W3(W3TO56), .W4(W4TO56), .W5(W5TO56), .W6(W6TO56), .W7(W7TO56), .W8(W8TO56), .W9(W9TO56), .W10(W10TO56), .W11(W11TO56), .W12(W12TO56), .W13(W13TO56), .W14(W14TO56), .W15(W15TO56), .W16(W16TO56), .W17(W17TO56), .W18(W18TO56), .W19(W19TO56), .W20(W20TO56), .W21(W21TO56), .W22(W22TO56), .W23(W23TO56), .W24(W24TO56), .W25(W25TO56), .W26(W26TO56), .W27(W27TO56), .W28(W28TO56), .W29(W29TO56), .W30(W30TO56), .W31(W31TO56), .W32(W32TO56), .W33(W33TO56), .W34(W34TO56), .W35(W35TO56), .W36(W36TO56), .W37(W37TO56), .W38(W38TO56), .W39(W39TO56), .W40(W40TO56), .W41(W41TO56), .W42(W42TO56), .W43(W43TO56), .W44(W44TO56), .W45(W45TO56), .W46(W46TO56), .W47(W47TO56), .W48(W48TO56), .W49(W49TO56), .W50(W50TO56), .W51(W51TO56), .W52(W52TO56), .W53(W53TO56), .W54(W54TO56), .W55(W55TO56), .W56(W56TO56), .W57(W57TO56), .W58(W58TO56), .W59(W59TO56), .W60(W60TO56), .W61(W61TO56), .W62(W62TO56), .W63(W63TO56), .W64(W64TO56)) neuron56(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out56));
neuron65in #(.BIAS(BIAS57), .W0(W0TO57), .W1(W1TO57), .W2(W2TO57), .W3(W3TO57), .W4(W4TO57), .W5(W5TO57), .W6(W6TO57), .W7(W7TO57), .W8(W8TO57), .W9(W9TO57), .W10(W10TO57), .W11(W11TO57), .W12(W12TO57), .W13(W13TO57), .W14(W14TO57), .W15(W15TO57), .W16(W16TO57), .W17(W17TO57), .W18(W18TO57), .W19(W19TO57), .W20(W20TO57), .W21(W21TO57), .W22(W22TO57), .W23(W23TO57), .W24(W24TO57), .W25(W25TO57), .W26(W26TO57), .W27(W27TO57), .W28(W28TO57), .W29(W29TO57), .W30(W30TO57), .W31(W31TO57), .W32(W32TO57), .W33(W33TO57), .W34(W34TO57), .W35(W35TO57), .W36(W36TO57), .W37(W37TO57), .W38(W38TO57), .W39(W39TO57), .W40(W40TO57), .W41(W41TO57), .W42(W42TO57), .W43(W43TO57), .W44(W44TO57), .W45(W45TO57), .W46(W46TO57), .W47(W47TO57), .W48(W48TO57), .W49(W49TO57), .W50(W50TO57), .W51(W51TO57), .W52(W52TO57), .W53(W53TO57), .W54(W54TO57), .W55(W55TO57), .W56(W56TO57), .W57(W57TO57), .W58(W58TO57), .W59(W59TO57), .W60(W60TO57), .W61(W61TO57), .W62(W62TO57), .W63(W63TO57), .W64(W64TO57)) neuron57(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out57));
neuron65in #(.BIAS(BIAS58), .W0(W0TO58), .W1(W1TO58), .W2(W2TO58), .W3(W3TO58), .W4(W4TO58), .W5(W5TO58), .W6(W6TO58), .W7(W7TO58), .W8(W8TO58), .W9(W9TO58), .W10(W10TO58), .W11(W11TO58), .W12(W12TO58), .W13(W13TO58), .W14(W14TO58), .W15(W15TO58), .W16(W16TO58), .W17(W17TO58), .W18(W18TO58), .W19(W19TO58), .W20(W20TO58), .W21(W21TO58), .W22(W22TO58), .W23(W23TO58), .W24(W24TO58), .W25(W25TO58), .W26(W26TO58), .W27(W27TO58), .W28(W28TO58), .W29(W29TO58), .W30(W30TO58), .W31(W31TO58), .W32(W32TO58), .W33(W33TO58), .W34(W34TO58), .W35(W35TO58), .W36(W36TO58), .W37(W37TO58), .W38(W38TO58), .W39(W39TO58), .W40(W40TO58), .W41(W41TO58), .W42(W42TO58), .W43(W43TO58), .W44(W44TO58), .W45(W45TO58), .W46(W46TO58), .W47(W47TO58), .W48(W48TO58), .W49(W49TO58), .W50(W50TO58), .W51(W51TO58), .W52(W52TO58), .W53(W53TO58), .W54(W54TO58), .W55(W55TO58), .W56(W56TO58), .W57(W57TO58), .W58(W58TO58), .W59(W59TO58), .W60(W60TO58), .W61(W61TO58), .W62(W62TO58), .W63(W63TO58), .W64(W64TO58)) neuron58(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out58));
neuron65in #(.BIAS(BIAS59), .W0(W0TO59), .W1(W1TO59), .W2(W2TO59), .W3(W3TO59), .W4(W4TO59), .W5(W5TO59), .W6(W6TO59), .W7(W7TO59), .W8(W8TO59), .W9(W9TO59), .W10(W10TO59), .W11(W11TO59), .W12(W12TO59), .W13(W13TO59), .W14(W14TO59), .W15(W15TO59), .W16(W16TO59), .W17(W17TO59), .W18(W18TO59), .W19(W19TO59), .W20(W20TO59), .W21(W21TO59), .W22(W22TO59), .W23(W23TO59), .W24(W24TO59), .W25(W25TO59), .W26(W26TO59), .W27(W27TO59), .W28(W28TO59), .W29(W29TO59), .W30(W30TO59), .W31(W31TO59), .W32(W32TO59), .W33(W33TO59), .W34(W34TO59), .W35(W35TO59), .W36(W36TO59), .W37(W37TO59), .W38(W38TO59), .W39(W39TO59), .W40(W40TO59), .W41(W41TO59), .W42(W42TO59), .W43(W43TO59), .W44(W44TO59), .W45(W45TO59), .W46(W46TO59), .W47(W47TO59), .W48(W48TO59), .W49(W49TO59), .W50(W50TO59), .W51(W51TO59), .W52(W52TO59), .W53(W53TO59), .W54(W54TO59), .W55(W55TO59), .W56(W56TO59), .W57(W57TO59), .W58(W58TO59), .W59(W59TO59), .W60(W60TO59), .W61(W61TO59), .W62(W62TO59), .W63(W63TO59), .W64(W64TO59)) neuron59(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out59));
neuron65in #(.BIAS(BIAS60), .W0(W0TO60), .W1(W1TO60), .W2(W2TO60), .W3(W3TO60), .W4(W4TO60), .W5(W5TO60), .W6(W6TO60), .W7(W7TO60), .W8(W8TO60), .W9(W9TO60), .W10(W10TO60), .W11(W11TO60), .W12(W12TO60), .W13(W13TO60), .W14(W14TO60), .W15(W15TO60), .W16(W16TO60), .W17(W17TO60), .W18(W18TO60), .W19(W19TO60), .W20(W20TO60), .W21(W21TO60), .W22(W22TO60), .W23(W23TO60), .W24(W24TO60), .W25(W25TO60), .W26(W26TO60), .W27(W27TO60), .W28(W28TO60), .W29(W29TO60), .W30(W30TO60), .W31(W31TO60), .W32(W32TO60), .W33(W33TO60), .W34(W34TO60), .W35(W35TO60), .W36(W36TO60), .W37(W37TO60), .W38(W38TO60), .W39(W39TO60), .W40(W40TO60), .W41(W41TO60), .W42(W42TO60), .W43(W43TO60), .W44(W44TO60), .W45(W45TO60), .W46(W46TO60), .W47(W47TO60), .W48(W48TO60), .W49(W49TO60), .W50(W50TO60), .W51(W51TO60), .W52(W52TO60), .W53(W53TO60), .W54(W54TO60), .W55(W55TO60), .W56(W56TO60), .W57(W57TO60), .W58(W58TO60), .W59(W59TO60), .W60(W60TO60), .W61(W61TO60), .W62(W62TO60), .W63(W63TO60), .W64(W64TO60)) neuron60(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out60));
neuron65in #(.BIAS(BIAS61), .W0(W0TO61), .W1(W1TO61), .W2(W2TO61), .W3(W3TO61), .W4(W4TO61), .W5(W5TO61), .W6(W6TO61), .W7(W7TO61), .W8(W8TO61), .W9(W9TO61), .W10(W10TO61), .W11(W11TO61), .W12(W12TO61), .W13(W13TO61), .W14(W14TO61), .W15(W15TO61), .W16(W16TO61), .W17(W17TO61), .W18(W18TO61), .W19(W19TO61), .W20(W20TO61), .W21(W21TO61), .W22(W22TO61), .W23(W23TO61), .W24(W24TO61), .W25(W25TO61), .W26(W26TO61), .W27(W27TO61), .W28(W28TO61), .W29(W29TO61), .W30(W30TO61), .W31(W31TO61), .W32(W32TO61), .W33(W33TO61), .W34(W34TO61), .W35(W35TO61), .W36(W36TO61), .W37(W37TO61), .W38(W38TO61), .W39(W39TO61), .W40(W40TO61), .W41(W41TO61), .W42(W42TO61), .W43(W43TO61), .W44(W44TO61), .W45(W45TO61), .W46(W46TO61), .W47(W47TO61), .W48(W48TO61), .W49(W49TO61), .W50(W50TO61), .W51(W51TO61), .W52(W52TO61), .W53(W53TO61), .W54(W54TO61), .W55(W55TO61), .W56(W56TO61), .W57(W57TO61), .W58(W58TO61), .W59(W59TO61), .W60(W60TO61), .W61(W61TO61), .W62(W62TO61), .W63(W63TO61), .W64(W64TO61)) neuron61(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out61));
neuron65in #(.BIAS(BIAS62), .W0(W0TO62), .W1(W1TO62), .W2(W2TO62), .W3(W3TO62), .W4(W4TO62), .W5(W5TO62), .W6(W6TO62), .W7(W7TO62), .W8(W8TO62), .W9(W9TO62), .W10(W10TO62), .W11(W11TO62), .W12(W12TO62), .W13(W13TO62), .W14(W14TO62), .W15(W15TO62), .W16(W16TO62), .W17(W17TO62), .W18(W18TO62), .W19(W19TO62), .W20(W20TO62), .W21(W21TO62), .W22(W22TO62), .W23(W23TO62), .W24(W24TO62), .W25(W25TO62), .W26(W26TO62), .W27(W27TO62), .W28(W28TO62), .W29(W29TO62), .W30(W30TO62), .W31(W31TO62), .W32(W32TO62), .W33(W33TO62), .W34(W34TO62), .W35(W35TO62), .W36(W36TO62), .W37(W37TO62), .W38(W38TO62), .W39(W39TO62), .W40(W40TO62), .W41(W41TO62), .W42(W42TO62), .W43(W43TO62), .W44(W44TO62), .W45(W45TO62), .W46(W46TO62), .W47(W47TO62), .W48(W48TO62), .W49(W49TO62), .W50(W50TO62), .W51(W51TO62), .W52(W52TO62), .W53(W53TO62), .W54(W54TO62), .W55(W55TO62), .W56(W56TO62), .W57(W57TO62), .W58(W58TO62), .W59(W59TO62), .W60(W60TO62), .W61(W61TO62), .W62(W62TO62), .W63(W63TO62), .W64(W64TO62)) neuron62(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out62));
neuron65in #(.BIAS(BIAS63), .W0(W0TO63), .W1(W1TO63), .W2(W2TO63), .W3(W3TO63), .W4(W4TO63), .W5(W5TO63), .W6(W6TO63), .W7(W7TO63), .W8(W8TO63), .W9(W9TO63), .W10(W10TO63), .W11(W11TO63), .W12(W12TO63), .W13(W13TO63), .W14(W14TO63), .W15(W15TO63), .W16(W16TO63), .W17(W17TO63), .W18(W18TO63), .W19(W19TO63), .W20(W20TO63), .W21(W21TO63), .W22(W22TO63), .W23(W23TO63), .W24(W24TO63), .W25(W25TO63), .W26(W26TO63), .W27(W27TO63), .W28(W28TO63), .W29(W29TO63), .W30(W30TO63), .W31(W31TO63), .W32(W32TO63), .W33(W33TO63), .W34(W34TO63), .W35(W35TO63), .W36(W36TO63), .W37(W37TO63), .W38(W38TO63), .W39(W39TO63), .W40(W40TO63), .W41(W41TO63), .W42(W42TO63), .W43(W43TO63), .W44(W44TO63), .W45(W45TO63), .W46(W46TO63), .W47(W47TO63), .W48(W48TO63), .W49(W49TO63), .W50(W50TO63), .W51(W51TO63), .W52(W52TO63), .W53(W53TO63), .W54(W54TO63), .W55(W55TO63), .W56(W56TO63), .W57(W57TO63), .W58(W58TO63), .W59(W59TO63), .W60(W60TO63), .W61(W61TO63), .W62(W62TO63), .W63(W63TO63), .W64(W64TO63)) neuron63(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out(out63));

endmodule

module layer64in1out(clk, rst, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, out0);

parameter signed BIAS0 = 0;
parameter signed W0TO0 = 0;
parameter signed W1TO0 = 0;
parameter signed W2TO0 = 0;
parameter signed W3TO0 = 0;
parameter signed W4TO0 = 0;
parameter signed W5TO0 = 0;
parameter signed W6TO0 = 0;
parameter signed W7TO0 = 0;
parameter signed W8TO0 = 0;
parameter signed W9TO0 = 0;
parameter signed W10TO0 = 0;
parameter signed W11TO0 = 0;
parameter signed W12TO0 = 0;
parameter signed W13TO0 = 0;
parameter signed W14TO0 = 0;
parameter signed W15TO0 = 0;
parameter signed W16TO0 = 0;
parameter signed W17TO0 = 0;
parameter signed W18TO0 = 0;
parameter signed W19TO0 = 0;
parameter signed W20TO0 = 0;
parameter signed W21TO0 = 0;
parameter signed W22TO0 = 0;
parameter signed W23TO0 = 0;
parameter signed W24TO0 = 0;
parameter signed W25TO0 = 0;
parameter signed W26TO0 = 0;
parameter signed W27TO0 = 0;
parameter signed W28TO0 = 0;
parameter signed W29TO0 = 0;
parameter signed W30TO0 = 0;
parameter signed W31TO0 = 0;
parameter signed W32TO0 = 0;
parameter signed W33TO0 = 0;
parameter signed W34TO0 = 0;
parameter signed W35TO0 = 0;
parameter signed W36TO0 = 0;
parameter signed W37TO0 = 0;
parameter signed W38TO0 = 0;
parameter signed W39TO0 = 0;
parameter signed W40TO0 = 0;
parameter signed W41TO0 = 0;
parameter signed W42TO0 = 0;
parameter signed W43TO0 = 0;
parameter signed W44TO0 = 0;
parameter signed W45TO0 = 0;
parameter signed W46TO0 = 0;
parameter signed W47TO0 = 0;
parameter signed W48TO0 = 0;
parameter signed W49TO0 = 0;
parameter signed W50TO0 = 0;
parameter signed W51TO0 = 0;
parameter signed W52TO0 = 0;
parameter signed W53TO0 = 0;
parameter signed W54TO0 = 0;
parameter signed W55TO0 = 0;
parameter signed W56TO0 = 0;
parameter signed W57TO0 = 0;
parameter signed W58TO0 = 0;
parameter signed W59TO0 = 0;
parameter signed W60TO0 = 0;
parameter signed W61TO0 = 0;
parameter signed W62TO0 = 0;
parameter signed W63TO0 = 0;

input wire clk;
input wire rst;

input signed [63:0] in0;
input signed [63:0] in1;
input signed [63:0] in2;
input signed [63:0] in3;
input signed [63:0] in4;
input signed [63:0] in5;
input signed [63:0] in6;
input signed [63:0] in7;
input signed [63:0] in8;
input signed [63:0] in9;
input signed [63:0] in10;
input signed [63:0] in11;
input signed [63:0] in12;
input signed [63:0] in13;
input signed [63:0] in14;
input signed [63:0] in15;
input signed [63:0] in16;
input signed [63:0] in17;
input signed [63:0] in18;
input signed [63:0] in19;
input signed [63:0] in20;
input signed [63:0] in21;
input signed [63:0] in22;
input signed [63:0] in23;
input signed [63:0] in24;
input signed [63:0] in25;
input signed [63:0] in26;
input signed [63:0] in27;
input signed [63:0] in28;
input signed [63:0] in29;
input signed [63:0] in30;
input signed [63:0] in31;
input signed [63:0] in32;
input signed [63:0] in33;
input signed [63:0] in34;
input signed [63:0] in35;
input signed [63:0] in36;
input signed [63:0] in37;
input signed [63:0] in38;
input signed [63:0] in39;
input signed [63:0] in40;
input signed [63:0] in41;
input signed [63:0] in42;
input signed [63:0] in43;
input signed [63:0] in44;
input signed [63:0] in45;
input signed [63:0] in46;
input signed [63:0] in47;
input signed [63:0] in48;
input signed [63:0] in49;
input signed [63:0] in50;
input signed [63:0] in51;
input signed [63:0] in52;
input signed [63:0] in53;
input signed [63:0] in54;
input signed [63:0] in55;
input signed [63:0] in56;
input signed [63:0] in57;
input signed [63:0] in58;
input signed [63:0] in59;
input signed [63:0] in60;
input signed [63:0] in61;
input signed [63:0] in62;
input signed [63:0] in63;

output signed [63:0] out0;

neuron64in #(.BIAS(BIAS0), .W0(W0TO0), .W1(W1TO0), .W2(W2TO0), .W3(W3TO0), .W4(W4TO0), .W5(W5TO0), .W6(W6TO0), .W7(W7TO0), .W8(W8TO0), .W9(W9TO0), .W10(W10TO0), .W11(W11TO0), .W12(W12TO0), .W13(W13TO0), .W14(W14TO0), .W15(W15TO0), .W16(W16TO0), .W17(W17TO0), .W18(W18TO0), .W19(W19TO0), .W20(W20TO0), .W21(W21TO0), .W22(W22TO0), .W23(W23TO0), .W24(W24TO0), .W25(W25TO0), .W26(W26TO0), .W27(W27TO0), .W28(W28TO0), .W29(W29TO0), .W30(W30TO0), .W31(W31TO0), .W32(W32TO0), .W33(W33TO0), .W34(W34TO0), .W35(W35TO0), .W36(W36TO0), .W37(W37TO0), .W38(W38TO0), .W39(W39TO0), .W40(W40TO0), .W41(W41TO0), .W42(W42TO0), .W43(W43TO0), .W44(W44TO0), .W45(W45TO0), .W46(W46TO0), .W47(W47TO0), .W48(W48TO0), .W49(W49TO0), .W50(W50TO0), .W51(W51TO0), .W52(W52TO0), .W53(W53TO0), .W54(W54TO0), .W55(W55TO0), .W56(W56TO0), .W57(W57TO0), .W58(W58TO0), .W59(W59TO0), .W60(W60TO0), .W61(W61TO0), .W62(W62TO0), .W63(W63TO0)) neuron0(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .out(out0));

endmodule

module network(clk, rst, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, out0);

input wire clk;
input wire rst;

input signed [63:0] in0;
input signed [63:0] in1;
input signed [63:0] in2;
input signed [63:0] in3;
input signed [63:0] in4;
input signed [63:0] in5;
input signed [63:0] in6;
input signed [63:0] in7;
input signed [63:0] in8;
input signed [63:0] in9;
input signed [63:0] in10;
input signed [63:0] in11;
input signed [63:0] in12;
input signed [63:0] in13;
input signed [63:0] in14;
input signed [63:0] in15;
input signed [63:0] in16;
input signed [63:0] in17;
input signed [63:0] in18;
input signed [63:0] in19;
input signed [63:0] in20;
input signed [63:0] in21;
input signed [63:0] in22;
input signed [63:0] in23;
input signed [63:0] in24;
input signed [63:0] in25;
input signed [63:0] in26;
input signed [63:0] in27;
input signed [63:0] in28;
input signed [63:0] in29;
input signed [63:0] in30;
input signed [63:0] in31;
input signed [63:0] in32;
input signed [63:0] in33;
input signed [63:0] in34;
input signed [63:0] in35;
input signed [63:0] in36;
input signed [63:0] in37;
input signed [63:0] in38;
input signed [63:0] in39;
input signed [63:0] in40;
input signed [63:0] in41;
input signed [63:0] in42;
input signed [63:0] in43;
input signed [63:0] in44;
input signed [63:0] in45;
input signed [63:0] in46;
input signed [63:0] in47;
input signed [63:0] in48;
input signed [63:0] in49;
input signed [63:0] in50;
input signed [63:0] in51;
input signed [63:0] in52;
input signed [63:0] in53;
input signed [63:0] in54;
input signed [63:0] in55;
input signed [63:0] in56;
input signed [63:0] in57;
input signed [63:0] in58;
input signed [63:0] in59;
input signed [63:0] in60;
input signed [63:0] in61;
input signed [63:0] in62;
input signed [63:0] in63;
input signed [63:0] in64;

output signed [63:0] out0;

wire[63:0] con0[0:63];

layer65in64out #(.BIAS0(-475950), .BIAS1(-682631), .BIAS2(-443746), .BIAS3(-81365), .BIAS4(-357998), .BIAS5(36786), .BIAS6(-476113), .BIAS7(952171), .BIAS8(465629), .BIAS9(-769451), .BIAS10(-227449), .BIAS11(257002), .BIAS12(-749883), .BIAS13(967097), .BIAS14(-113549), .BIAS15(579117), .BIAS16(588237), .BIAS17(-277476), .BIAS18(-167791), .BIAS19(168516), .BIAS20(520344), .BIAS21(-624382), .BIAS22(-423665), .BIAS23(340438), .BIAS24(-702), .BIAS25(-642862), .BIAS26(-173716), .BIAS27(-601609), .BIAS28(63399), .BIAS29(664741), .BIAS30(-629497), .BIAS31(914718), .BIAS32(-149170), .BIAS33(8014), .BIAS34(20942), .BIAS35(-968416), .BIAS36(463380), .BIAS37(986610), .BIAS38(-674244), .BIAS39(-746729), .BIAS40(-250331), .BIAS41(386439), .BIAS42(-994197), .BIAS43(-261541), .BIAS44(-882640), .BIAS45(578672), .BIAS46(-300461), .BIAS47(405047), .BIAS48(-17541), .BIAS49(945745), .BIAS50(671936), .BIAS51(220475), .BIAS52(129038), .BIAS53(994778), .BIAS54(-490551), .BIAS55(-971243), .BIAS56(-821909), .BIAS57(877965), .BIAS58(946919), .BIAS59(-17036), .BIAS60(-318127), .BIAS61(445715), .BIAS62(-978205), .BIAS63(519906), .W0TO0(342806), .W0TO1(-619108), .W0TO2(332929), .W0TO3(822245), .W0TO4(-675764), .W0TO5(821157), .W0TO6(-351283), .W0TO7(400597), .W0TO8(-469098), .W0TO9(37917), .W0TO10(-645063), .W0TO11(-64307), .W0TO12(-102070), .W0TO13(-207870), .W0TO14(583851), .W0TO15(-13203), .W0TO16(447896), .W0TO17(586046), .W0TO18(-296951), .W0TO19(819307), .W0TO20(425775), .W0TO21(794495), .W0TO22(-159582), .W0TO23(-64967), .W0TO24(807854), .W0TO25(267097), .W0TO26(65659), .W0TO27(-524977), .W0TO28(893008), .W0TO29(118860), .W0TO30(514703), .W0TO31(-527701), .W0TO32(-140482), .W0TO33(-211772), .W0TO34(21419), .W0TO35(-749193), .W0TO36(367306), .W0TO37(-944620), .W0TO38(-532313), .W0TO39(472884), .W0TO40(868420), .W0TO41(227208), .W0TO42(-185043), .W0TO43(707833), .W0TO44(985664), .W0TO45(-409259), .W0TO46(-219664), .W0TO47(397914), .W0TO48(-285960), .W0TO49(-936149), .W0TO50(-301716), .W0TO51(-30481), .W0TO52(-903529), .W0TO53(830051), .W0TO54(451133), .W0TO55(544923), .W0TO56(-807099), .W0TO57(-925539), .W0TO58(-480374), .W0TO59(-748984), .W0TO60(-523700), .W0TO61(364347), .W0TO62(-37562), .W0TO63(873017), .W1TO0(162797), .W1TO1(-627784), .W1TO2(-626143), .W1TO3(-322892), .W1TO4(-134464), .W1TO5(-846458), .W1TO6(272017), .W1TO7(-883180), .W1TO8(447360), .W1TO9(320204), .W1TO10(-982362), .W1TO11(526363), .W1TO12(-322735), .W1TO13(552426), .W1TO14(-328406), .W1TO15(161084), .W1TO16(-656045), .W1TO17(692435), .W1TO18(-458193), .W1TO19(489278), .W1TO20(126839), .W1TO21(800176), .W1TO22(96644), .W1TO23(-949716), .W1TO24(-838720), .W1TO25(911118), .W1TO26(-87936), .W1TO27(-705305), .W1TO28(349922), .W1TO29(247333), .W1TO30(100412), .W1TO31(811501), .W1TO32(796638), .W1TO33(-475194), .W1TO34(438314), .W1TO35(-29706), .W1TO36(-438229), .W1TO37(-883440), .W1TO38(-589882), .W1TO39(280078), .W1TO40(-428050), .W1TO41(-114922), .W1TO42(-308108), .W1TO43(-525), .W1TO44(310144), .W1TO45(898830), .W1TO46(-933851), .W1TO47(112678), .W1TO48(281600), .W1TO49(-683117), .W1TO50(452895), .W1TO51(-242959), .W1TO52(23106), .W1TO53(156482), .W1TO54(690562), .W1TO55(403658), .W1TO56(258379), .W1TO57(-897313), .W1TO58(-908179), .W1TO59(58030), .W1TO60(566086), .W1TO61(406156), .W1TO62(-606761), .W1TO63(-456510), .W2TO0(-569498), .W2TO1(-183305), .W2TO2(310552), .W2TO3(-459359), .W2TO4(-439110), .W2TO5(563540), .W2TO6(704233), .W2TO7(94872), .W2TO8(448229), .W2TO9(-133663), .W2TO10(641067), .W2TO11(648659), .W2TO12(-966916), .W2TO13(466080), .W2TO14(434486), .W2TO15(438515), .W2TO16(572146), .W2TO17(874383), .W2TO18(316326), .W2TO19(-625003), .W2TO20(376411), .W2TO21(980782), .W2TO22(828741), .W2TO23(730164), .W2TO24(-906593), .W2TO25(-984321), .W2TO26(499013), .W2TO27(467080), .W2TO28(416740), .W2TO29(-685834), .W2TO30(-762907), .W2TO31(-679195), .W2TO32(646346), .W2TO33(-192563), .W2TO34(-641738), .W2TO35(262913), .W2TO36(-923755), .W2TO37(-811793), .W2TO38(-776623), .W2TO39(378906), .W2TO40(234532), .W2TO41(147606), .W2TO42(652219), .W2TO43(489556), .W2TO44(-546697), .W2TO45(-824222), .W2TO46(1872), .W2TO47(-372615), .W2TO48(-464052), .W2TO49(18884), .W2TO50(403257), .W2TO51(814368), .W2TO52(-92413), .W2TO53(66417), .W2TO54(617630), .W2TO55(-221549), .W2TO56(485964), .W2TO57(969821), .W2TO58(-578514), .W2TO59(156830), .W2TO60(441435), .W2TO61(-732872), .W2TO62(626018), .W2TO63(474231), .W3TO0(488797), .W3TO1(687080), .W3TO2(499518), .W3TO3(482228), .W3TO4(283811), .W3TO5(279448), .W3TO6(655705), .W3TO7(668063), .W3TO8(-557017), .W3TO9(324351), .W3TO10(-641559), .W3TO11(643094), .W3TO12(-936338), .W3TO13(-931506), .W3TO14(-961140), .W3TO15(291161), .W3TO16(63311), .W3TO17(-944877), .W3TO18(-947114), .W3TO19(495364), .W3TO20(497392), .W3TO21(-537157), .W3TO22(569056), .W3TO23(688476), .W3TO24(660946), .W3TO25(110206), .W3TO26(383608), .W3TO27(544159), .W3TO28(477489), .W3TO29(-185860), .W3TO30(342669), .W3TO31(393854), .W3TO32(630127), .W3TO33(-301341), .W3TO34(47453), .W3TO35(-616405), .W3TO36(-495109), .W3TO37(82925), .W3TO38(-397002), .W3TO39(290047), .W3TO40(-902195), .W3TO41(-781243), .W3TO42(515355), .W3TO43(-114294), .W3TO44(939408), .W3TO45(-754929), .W3TO46(-284352), .W3TO47(846991), .W3TO48(671750), .W3TO49(956329), .W3TO50(-608918), .W3TO51(-281283), .W3TO52(290461), .W3TO53(-445858), .W3TO54(-906232), .W3TO55(163124), .W3TO56(-624702), .W3TO57(578663), .W3TO58(-239300), .W3TO59(-347074), .W3TO60(302607), .W3TO61(249562), .W3TO62(-376847), .W3TO63(495852), .W4TO0(-193618), .W4TO1(529930), .W4TO2(-911563), .W4TO3(819696), .W4TO4(292726), .W4TO5(-94735), .W4TO6(-955909), .W4TO7(-582360), .W4TO8(226582), .W4TO9(856112), .W4TO10(208498), .W4TO11(122887), .W4TO12(-171351), .W4TO13(671747), .W4TO14(162547), .W4TO15(489237), .W4TO16(-508481), .W4TO17(-771181), .W4TO18(979556), .W4TO19(-934831), .W4TO20(-557033), .W4TO21(-169434), .W4TO22(-521461), .W4TO23(-469027), .W4TO24(111522), .W4TO25(219903), .W4TO26(213508), .W4TO27(522914), .W4TO28(-569438), .W4TO29(787144), .W4TO30(320745), .W4TO31(-909517), .W4TO32(193768), .W4TO33(-245237), .W4TO34(-311394), .W4TO35(-602477), .W4TO36(430838), .W4TO37(954595), .W4TO38(-444286), .W4TO39(310988), .W4TO40(-125524), .W4TO41(-133716), .W4TO42(-788508), .W4TO43(-496998), .W4TO44(736331), .W4TO45(-768251), .W4TO46(-366882), .W4TO47(429761), .W4TO48(-241126), .W4TO49(-459091), .W4TO50(893807), .W4TO51(820019), .W4TO52(220537), .W4TO53(992332), .W4TO54(973199), .W4TO55(755911), .W4TO56(2952), .W4TO57(623305), .W4TO58(591806), .W4TO59(-644827), .W4TO60(214825), .W4TO61(-804243), .W4TO62(-542357), .W4TO63(-713515), .W5TO0(-380865), .W5TO1(-93135), .W5TO2(-407236), .W5TO3(119017), .W5TO4(743574), .W5TO5(-585844), .W5TO6(-884797), .W5TO7(816115), .W5TO8(-319686), .W5TO9(682500), .W5TO10(864670), .W5TO11(619015), .W5TO12(-874487), .W5TO13(-194302), .W5TO14(-486483), .W5TO15(288189), .W5TO16(145566), .W5TO17(851148), .W5TO18(-212242), .W5TO19(675284), .W5TO20(364310), .W5TO21(-332569), .W5TO22(-431875), .W5TO23(410414), .W5TO24(142611), .W5TO25(942637), .W5TO26(-560527), .W5TO27(-528056), .W5TO28(387479), .W5TO29(322880), .W5TO30(839730), .W5TO31(843951), .W5TO32(-493694), .W5TO33(74939), .W5TO34(-208935), .W5TO35(-816847), .W5TO36(-453814), .W5TO37(-828115), .W5TO38(952633), .W5TO39(799714), .W5TO40(667608), .W5TO41(958833), .W5TO42(194857), .W5TO43(359679), .W5TO44(-556738), .W5TO45(852083), .W5TO46(-922955), .W5TO47(264264), .W5TO48(-920587), .W5TO49(946731), .W5TO50(751200), .W5TO51(7473), .W5TO52(178748), .W5TO53(-438348), .W5TO54(-693769), .W5TO55(658651), .W5TO56(-737319), .W5TO57(-735573), .W5TO58(-311437), .W5TO59(976316), .W5TO60(-33431), .W5TO61(-384964), .W5TO62(-499838), .W5TO63(563030), .W6TO0(-707607), .W6TO1(-123101), .W6TO2(736147), .W6TO3(-972179), .W6TO4(514866), .W6TO5(958001), .W6TO6(-533882), .W6TO7(481329), .W6TO8(600592), .W6TO9(742440), .W6TO10(392095), .W6TO11(-557959), .W6TO12(-837286), .W6TO13(118282), .W6TO14(118806), .W6TO15(-200689), .W6TO16(91942), .W6TO17(-667268), .W6TO18(-653229), .W6TO19(429567), .W6TO20(993580), .W6TO21(601960), .W6TO22(-667788), .W6TO23(547850), .W6TO24(-419168), .W6TO25(854987), .W6TO26(-53949), .W6TO27(-203955), .W6TO28(-800900), .W6TO29(10083), .W6TO30(-823906), .W6TO31(369488), .W6TO32(-724597), .W6TO33(-59870), .W6TO34(-504969), .W6TO35(998995), .W6TO36(-455024), .W6TO37(170333), .W6TO38(-971190), .W6TO39(222200), .W6TO40(21856), .W6TO41(-34400), .W6TO42(-194311), .W6TO43(778198), .W6TO44(-633390), .W6TO45(387182), .W6TO46(555221), .W6TO47(468733), .W6TO48(213905), .W6TO49(400809), .W6TO50(-518512), .W6TO51(-829741), .W6TO52(820746), .W6TO53(71270), .W6TO54(-517468), .W6TO55(687157), .W6TO56(632164), .W6TO57(-522998), .W6TO58(744244), .W6TO59(-347212), .W6TO60(-235808), .W6TO61(-190064), .W6TO62(12324), .W6TO63(-519048), .W7TO0(-52285), .W7TO1(-476489), .W7TO2(-217707), .W7TO3(775401), .W7TO4(-313942), .W7TO5(-713949), .W7TO6(451188), .W7TO7(-424809), .W7TO8(546707), .W7TO9(993886), .W7TO10(116118), .W7TO11(-654657), .W7TO12(-129902), .W7TO13(-176177), .W7TO14(-969422), .W7TO15(-846021), .W7TO16(376484), .W7TO17(99333), .W7TO18(864911), .W7TO19(189480), .W7TO20(380113), .W7TO21(75947), .W7TO22(155946), .W7TO23(-922537), .W7TO24(-489675), .W7TO25(220283), .W7TO26(-856977), .W7TO27(-93002), .W7TO28(484116), .W7TO29(-943143), .W7TO30(757503), .W7TO31(479796), .W7TO32(257276), .W7TO33(-417011), .W7TO34(-289206), .W7TO35(-716116), .W7TO36(-487307), .W7TO37(348012), .W7TO38(-946327), .W7TO39(868728), .W7TO40(-832941), .W7TO41(-945425), .W7TO42(-708794), .W7TO43(753278), .W7TO44(-615784), .W7TO45(-457647), .W7TO46(-115807), .W7TO47(-870453), .W7TO48(579868), .W7TO49(-380370), .W7TO50(590676), .W7TO51(-236346), .W7TO52(-858694), .W7TO53(645193), .W7TO54(342964), .W7TO55(49143), .W7TO56(-518151), .W7TO57(892866), .W7TO58(-36918), .W7TO59(835412), .W7TO60(588665), .W7TO61(355096), .W7TO62(34469), .W7TO63(959269), .W8TO0(-880591), .W8TO1(740893), .W8TO2(-905220), .W8TO3(-206954), .W8TO4(142965), .W8TO5(-28665), .W8TO6(-142754), .W8TO7(-123669), .W8TO8(-776742), .W8TO9(-721495), .W8TO10(-395752), .W8TO11(783883), .W8TO12(560771), .W8TO13(-568191), .W8TO14(-814734), .W8TO15(38394), .W8TO16(-644268), .W8TO17(-382548), .W8TO18(-664004), .W8TO19(-305819), .W8TO20(219865), .W8TO21(949829), .W8TO22(333481), .W8TO23(-183649), .W8TO24(-303174), .W8TO25(-275556), .W8TO26(801927), .W8TO27(-319809), .W8TO28(-872611), .W8TO29(2071), .W8TO30(-827066), .W8TO31(-835765), .W8TO32(925325), .W8TO33(-83864), .W8TO34(881090), .W8TO35(477225), .W8TO36(281495), .W8TO37(-80832), .W8TO38(-843074), .W8TO39(427622), .W8TO40(-397193), .W8TO41(548914), .W8TO42(-386076), .W8TO43(-12605), .W8TO44(261176), .W8TO45(-657663), .W8TO46(254925), .W8TO47(-776350), .W8TO48(-290679), .W8TO49(-197319), .W8TO50(-524413), .W8TO51(966429), .W8TO52(-877148), .W8TO53(778198), .W8TO54(269344), .W8TO55(920970), .W8TO56(164421), .W8TO57(421497), .W8TO58(712088), .W8TO59(604675), .W8TO60(-607924), .W8TO61(38474), .W8TO62(-330275), .W8TO63(878821), .W9TO0(290190), .W9TO1(37641), .W9TO2(325620), .W9TO3(-746657), .W9TO4(698502), .W9TO5(-378362), .W9TO6(-830619), .W9TO7(-440703), .W9TO8(252556), .W9TO9(-474516), .W9TO10(-853280), .W9TO11(933522), .W9TO12(349422), .W9TO13(-696669), .W9TO14(293065), .W9TO15(-769188), .W9TO16(-670988), .W9TO17(-764079), .W9TO18(-177383), .W9TO19(946025), .W9TO20(-729305), .W9TO21(-744141), .W9TO22(-666208), .W9TO23(267784), .W9TO24(375647), .W9TO25(235548), .W9TO26(-947053), .W9TO27(176352), .W9TO28(-911039), .W9TO29(274031), .W9TO30(-314919), .W9TO31(922737), .W9TO32(752910), .W9TO33(510239), .W9TO34(658372), .W9TO35(49947), .W9TO36(-192274), .W9TO37(-785566), .W9TO38(-4124), .W9TO39(-637069), .W9TO40(568408), .W9TO41(-703696), .W9TO42(-754760), .W9TO43(691538), .W9TO44(878175), .W9TO45(-100614), .W9TO46(-701895), .W9TO47(96547), .W9TO48(-695917), .W9TO49(-388490), .W9TO50(866460), .W9TO51(-863045), .W9TO52(-902325), .W9TO53(-779044), .W9TO54(-74802), .W9TO55(-584275), .W9TO56(814700), .W9TO57(-291364), .W9TO58(-220277), .W9TO59(-384551), .W9TO60(165747), .W9TO61(748671), .W9TO62(-699294), .W9TO63(431360), .W10TO0(527558), .W10TO1(476459), .W10TO2(-676241), .W10TO3(131815), .W10TO4(183460), .W10TO5(-897290), .W10TO6(-22043), .W10TO7(500854), .W10TO8(-913579), .W10TO9(177425), .W10TO10(209966), .W10TO11(-577619), .W10TO12(-853186), .W10TO13(292392), .W10TO14(568899), .W10TO15(150529), .W10TO16(-518450), .W10TO17(-639192), .W10TO18(-714956), .W10TO19(1139), .W10TO20(-771637), .W10TO21(-874705), .W10TO22(-756749), .W10TO23(-823163), .W10TO24(321920), .W10TO25(-183063), .W10TO26(293871), .W10TO27(-277883), .W10TO28(427596), .W10TO29(-6009), .W10TO30(582270), .W10TO31(916939), .W10TO32(-542999), .W10TO33(-550300), .W10TO34(73957), .W10TO35(-353583), .W10TO36(531762), .W10TO37(636640), .W10TO38(-69239), .W10TO39(-905165), .W10TO40(759493), .W10TO41(779108), .W10TO42(892432), .W10TO43(621814), .W10TO44(798473), .W10TO45(900265), .W10TO46(754777), .W10TO47(920299), .W10TO48(-105905), .W10TO49(680264), .W10TO50(-493573), .W10TO51(551204), .W10TO52(848461), .W10TO53(-293942), .W10TO54(-381808), .W10TO55(466820), .W10TO56(540829), .W10TO57(-65715), .W10TO58(230706), .W10TO59(348641), .W10TO60(-982270), .W10TO61(-261719), .W10TO62(-487733), .W10TO63(686309), .W11TO0(-558703), .W11TO1(963149), .W11TO2(992062), .W11TO3(206609), .W11TO4(-627645), .W11TO5(66269), .W11TO6(979595), .W11TO7(-282970), .W11TO8(-650713), .W11TO9(718362), .W11TO10(623164), .W11TO11(-998337), .W11TO12(-228861), .W11TO13(563075), .W11TO14(-84334), .W11TO15(377903), .W11TO16(714432), .W11TO17(245277), .W11TO18(528631), .W11TO19(265838), .W11TO20(-925030), .W11TO21(-515597), .W11TO22(404481), .W11TO23(-801729), .W11TO24(592498), .W11TO25(-648173), .W11TO26(-971714), .W11TO27(26585), .W11TO28(56369), .W11TO29(-39641), .W11TO30(-500939), .W11TO31(-736746), .W11TO32(-122334), .W11TO33(-671451), .W11TO34(-986149), .W11TO35(830145), .W11TO36(-170101), .W11TO37(813913), .W11TO38(147423), .W11TO39(-278955), .W11TO40(230153), .W11TO41(754369), .W11TO42(-643968), .W11TO43(-506159), .W11TO44(-51722), .W11TO45(-554393), .W11TO46(-6731), .W11TO47(-176373), .W11TO48(-329270), .W11TO49(-227179), .W11TO50(990217), .W11TO51(-5427), .W11TO52(-910688), .W11TO53(996558), .W11TO54(625089), .W11TO55(-352536), .W11TO56(-153813), .W11TO57(476723), .W11TO58(-310601), .W11TO59(-152348), .W11TO60(-299652), .W11TO61(-80285), .W11TO62(61592), .W11TO63(895622), .W12TO0(-433249), .W12TO1(499214), .W12TO2(-682491), .W12TO3(-737085), .W12TO4(-151087), .W12TO5(665833), .W12TO6(-364119), .W12TO7(734144), .W12TO8(-598252), .W12TO9(-332632), .W12TO10(170296), .W12TO11(488030), .W12TO12(344929), .W12TO13(-490942), .W12TO14(454857), .W12TO15(-411277), .W12TO16(-546496), .W12TO17(-801659), .W12TO18(-292432), .W12TO19(741566), .W12TO20(587970), .W12TO21(-632798), .W12TO22(-468971), .W12TO23(402380), .W12TO24(963291), .W12TO25(184493), .W12TO26(-420787), .W12TO27(-938741), .W12TO28(-57598), .W12TO29(-858639), .W12TO30(-711040), .W12TO31(666322), .W12TO32(758890), .W12TO33(376122), .W12TO34(-975185), .W12TO35(-352967), .W12TO36(832052), .W12TO37(973679), .W12TO38(312562), .W12TO39(592690), .W12TO40(119254), .W12TO41(-89015), .W12TO42(-198246), .W12TO43(273695), .W12TO44(-897167), .W12TO45(197976), .W12TO46(556695), .W12TO47(-696303), .W12TO48(-315518), .W12TO49(-835301), .W12TO50(-865200), .W12TO51(-534087), .W12TO52(-945771), .W12TO53(635677), .W12TO54(354349), .W12TO55(324388), .W12TO56(933994), .W12TO57(-57458), .W12TO58(314372), .W12TO59(532043), .W12TO60(-742375), .W12TO61(373658), .W12TO62(468349), .W12TO63(79586), .W13TO0(812851), .W13TO1(-41904), .W13TO2(700036), .W13TO3(689413), .W13TO4(699357), .W13TO5(823875), .W13TO6(459519), .W13TO7(691149), .W13TO8(-254011), .W13TO9(-114592), .W13TO10(502064), .W13TO11(-391772), .W13TO12(-208114), .W13TO13(-575794), .W13TO14(-171361), .W13TO15(-419160), .W13TO16(109721), .W13TO17(-197077), .W13TO18(-741655), .W13TO19(-968737), .W13TO20(726680), .W13TO21(-500570), .W13TO22(-106529), .W13TO23(-370444), .W13TO24(-778109), .W13TO25(934034), .W13TO26(-27653), .W13TO27(569982), .W13TO28(-414533), .W13TO29(-414421), .W13TO30(-694185), .W13TO31(-400065), .W13TO32(-711318), .W13TO33(940197), .W13TO34(703407), .W13TO35(-251487), .W13TO36(614215), .W13TO37(773543), .W13TO38(-994234), .W13TO39(1454), .W13TO40(-898232), .W13TO41(-96525), .W13TO42(620602), .W13TO43(417985), .W13TO44(364447), .W13TO45(386589), .W13TO46(606199), .W13TO47(497441), .W13TO48(-58860), .W13TO49(533580), .W13TO50(-327426), .W13TO51(-771654), .W13TO52(45225), .W13TO53(453578), .W13TO54(687656), .W13TO55(-990110), .W13TO56(-958191), .W13TO57(-142530), .W13TO58(-536353), .W13TO59(-288868), .W13TO60(-813280), .W13TO61(448403), .W13TO62(-767619), .W13TO63(41320), .W14TO0(939166), .W14TO1(720376), .W14TO2(-821481), .W14TO3(-866485), .W14TO4(155287), .W14TO5(-23195), .W14TO6(-416875), .W14TO7(-225900), .W14TO8(826647), .W14TO9(-616931), .W14TO10(743542), .W14TO11(882262), .W14TO12(810671), .W14TO13(-271915), .W14TO14(-289348), .W14TO15(854792), .W14TO16(840491), .W14TO17(-317613), .W14TO18(-681181), .W14TO19(357970), .W14TO20(-130270), .W14TO21(65804), .W14TO22(310371), .W14TO23(896441), .W14TO24(-47903), .W14TO25(-149042), .W14TO26(-494422), .W14TO27(-68548), .W14TO28(131588), .W14TO29(27853), .W14TO30(-735246), .W14TO31(759589), .W14TO32(-341395), .W14TO33(-996757), .W14TO34(-201116), .W14TO35(-852155), .W14TO36(-917184), .W14TO37(-166960), .W14TO38(496538), .W14TO39(603976), .W14TO40(245822), .W14TO41(-606873), .W14TO42(-283398), .W14TO43(194193), .W14TO44(914128), .W14TO45(651416), .W14TO46(842483), .W14TO47(-40603), .W14TO48(-653877), .W14TO49(-995447), .W14TO50(-206076), .W14TO51(112879), .W14TO52(651389), .W14TO53(-962603), .W14TO54(573265), .W14TO55(-331947), .W14TO56(402289), .W14TO57(160786), .W14TO58(996465), .W14TO59(-306664), .W14TO60(543071), .W14TO61(-570482), .W14TO62(597783), .W14TO63(-23022), .W15TO0(-467740), .W15TO1(-838479), .W15TO2(800385), .W15TO3(573962), .W15TO4(773285), .W15TO5(-573805), .W15TO6(-476), .W15TO7(-881130), .W15TO8(-736009), .W15TO9(838668), .W15TO10(230040), .W15TO11(46412), .W15TO12(-510730), .W15TO13(280022), .W15TO14(-846897), .W15TO15(-132658), .W15TO16(-558487), .W15TO17(264708), .W15TO18(107684), .W15TO19(965295), .W15TO20(69137), .W15TO21(634697), .W15TO22(691387), .W15TO23(691891), .W15TO24(182731), .W15TO25(648505), .W15TO26(432237), .W15TO27(283647), .W15TO28(434573), .W15TO29(-538417), .W15TO30(969800), .W15TO31(-520273), .W15TO32(507259), .W15TO33(691406), .W15TO34(185597), .W15TO35(308486), .W15TO36(432146), .W15TO37(139697), .W15TO38(671132), .W15TO39(964755), .W15TO40(471519), .W15TO41(-185739), .W15TO42(245327), .W15TO43(-928293), .W15TO44(111989), .W15TO45(-30458), .W15TO46(-862099), .W15TO47(-524600), .W15TO48(-366420), .W15TO49(588503), .W15TO50(-948998), .W15TO51(890245), .W15TO52(367750), .W15TO53(-422432), .W15TO54(-739228), .W15TO55(188723), .W15TO56(482638), .W15TO57(168978), .W15TO58(-790651), .W15TO59(971021), .W15TO60(76274), .W15TO61(-437635), .W15TO62(234247), .W15TO63(-874125), .W16TO0(-934626), .W16TO1(608126), .W16TO2(-475800), .W16TO3(896109), .W16TO4(-869966), .W16TO5(-74571), .W16TO6(-480710), .W16TO7(275262), .W16TO8(160526), .W16TO9(-216539), .W16TO10(47673), .W16TO11(-692677), .W16TO12(-522991), .W16TO13(730687), .W16TO14(722982), .W16TO15(974408), .W16TO16(-124483), .W16TO17(-869462), .W16TO18(-350475), .W16TO19(-828288), .W16TO20(562606), .W16TO21(650662), .W16TO22(-938746), .W16TO23(328502), .W16TO24(404408), .W16TO25(-522246), .W16TO26(-120831), .W16TO27(996568), .W16TO28(751420), .W16TO29(353364), .W16TO30(270896), .W16TO31(688603), .W16TO32(-265288), .W16TO33(-180321), .W16TO34(890504), .W16TO35(-81654), .W16TO36(-326351), .W16TO37(344748), .W16TO38(-118852), .W16TO39(506454), .W16TO40(-217983), .W16TO41(210587), .W16TO42(-619756), .W16TO43(-736738), .W16TO44(767855), .W16TO45(985101), .W16TO46(-499424), .W16TO47(-371640), .W16TO48(-397473), .W16TO49(366469), .W16TO50(-670693), .W16TO51(437216), .W16TO52(202555), .W16TO53(-796970), .W16TO54(201078), .W16TO55(537010), .W16TO56(-879890), .W16TO57(-862722), .W16TO58(993768), .W16TO59(345268), .W16TO60(-927717), .W16TO61(-108232), .W16TO62(90424), .W16TO63(-158753), .W17TO0(250982), .W17TO1(642268), .W17TO2(-210027), .W17TO3(-500471), .W17TO4(36483), .W17TO5(-986609), .W17TO6(-590214), .W17TO7(319942), .W17TO8(-425832), .W17TO9(-446537), .W17TO10(145291), .W17TO11(-132123), .W17TO12(-711743), .W17TO13(989978), .W17TO14(937186), .W17TO15(-56834), .W17TO16(480475), .W17TO17(324081), .W17TO18(430778), .W17TO19(34433), .W17TO20(-506453), .W17TO21(6562), .W17TO22(910851), .W17TO23(423169), .W17TO24(-983535), .W17TO25(-181801), .W17TO26(-129552), .W17TO27(754172), .W17TO28(-143127), .W17TO29(-355828), .W17TO30(541864), .W17TO31(838512), .W17TO32(-695696), .W17TO33(994940), .W17TO34(846039), .W17TO35(-335556), .W17TO36(18728), .W17TO37(-743731), .W17TO38(839937), .W17TO39(-152281), .W17TO40(-540079), .W17TO41(-579784), .W17TO42(149696), .W17TO43(755817), .W17TO44(-246274), .W17TO45(262375), .W17TO46(697394), .W17TO47(-953925), .W17TO48(594414), .W17TO49(700907), .W17TO50(-476518), .W17TO51(-560860), .W17TO52(161321), .W17TO53(172169), .W17TO54(-599021), .W17TO55(-68290), .W17TO56(108173), .W17TO57(-635565), .W17TO58(-352234), .W17TO59(212822), .W17TO60(-653476), .W17TO61(-115301), .W17TO62(-108800), .W17TO63(838605), .W18TO0(444477), .W18TO1(365501), .W18TO2(-490351), .W18TO3(363890), .W18TO4(-981680), .W18TO5(-156998), .W18TO6(955441), .W18TO7(-344280), .W18TO8(868630), .W18TO9(540265), .W18TO10(-443385), .W18TO11(-519721), .W18TO12(-696545), .W18TO13(47145), .W18TO14(45986), .W18TO15(-184104), .W18TO16(646056), .W18TO17(655915), .W18TO18(63234), .W18TO19(381280), .W18TO20(-14093), .W18TO21(-39953), .W18TO22(232865), .W18TO23(-565935), .W18TO24(-738799), .W18TO25(124036), .W18TO26(-377668), .W18TO27(-18803), .W18TO28(-416143), .W18TO29(-470348), .W18TO30(-155431), .W18TO31(-995853), .W18TO32(-458513), .W18TO33(-263164), .W18TO34(-17687), .W18TO35(891916), .W18TO36(111775), .W18TO37(720358), .W18TO38(194805), .W18TO39(-186487), .W18TO40(-965242), .W18TO41(859088), .W18TO42(-280283), .W18TO43(806410), .W18TO44(655427), .W18TO45(-855011), .W18TO46(-739098), .W18TO47(-433601), .W18TO48(-82153), .W18TO49(286470), .W18TO50(777815), .W18TO51(-142093), .W18TO52(486842), .W18TO53(827249), .W18TO54(-733773), .W18TO55(885607), .W18TO56(592875), .W18TO57(491043), .W18TO58(-108049), .W18TO59(-851778), .W18TO60(-479678), .W18TO61(319995), .W18TO62(-951761), .W18TO63(542726), .W19TO0(946285), .W19TO1(-754049), .W19TO2(290155), .W19TO3(698266), .W19TO4(408300), .W19TO5(691494), .W19TO6(865169), .W19TO7(616730), .W19TO8(-98488), .W19TO9(167415), .W19TO10(-24655), .W19TO11(227300), .W19TO12(29186), .W19TO13(280051), .W19TO14(594545), .W19TO15(909994), .W19TO16(5223), .W19TO17(-102147), .W19TO18(-527588), .W19TO19(800884), .W19TO20(603176), .W19TO21(-244405), .W19TO22(-624721), .W19TO23(-110260), .W19TO24(880120), .W19TO25(-247961), .W19TO26(-359758), .W19TO27(775750), .W19TO28(792621), .W19TO29(-251008), .W19TO30(899391), .W19TO31(676006), .W19TO32(174784), .W19TO33(-508644), .W19TO34(-527304), .W19TO35(-341411), .W19TO36(961840), .W19TO37(120801), .W19TO38(540173), .W19TO39(-100806), .W19TO40(731703), .W19TO41(907244), .W19TO42(390180), .W19TO43(40162), .W19TO44(-622781), .W19TO45(630129), .W19TO46(688181), .W19TO47(887547), .W19TO48(727519), .W19TO49(-184975), .W19TO50(-396862), .W19TO51(-51571), .W19TO52(953488), .W19TO53(661721), .W19TO54(-744145), .W19TO55(672817), .W19TO56(-210466), .W19TO57(953126), .W19TO58(998669), .W19TO59(462740), .W19TO60(679127), .W19TO61(-572770), .W19TO62(-288876), .W19TO63(689729), .W20TO0(-363425), .W20TO1(-10648), .W20TO2(530034), .W20TO3(-116625), .W20TO4(145124), .W20TO5(126494), .W20TO6(757906), .W20TO7(582780), .W20TO8(515699), .W20TO9(-344067), .W20TO10(-57209), .W20TO11(909286), .W20TO12(-720117), .W20TO13(378319), .W20TO14(-614957), .W20TO15(-473956), .W20TO16(-154216), .W20TO17(-496191), .W20TO18(-29627), .W20TO19(425920), .W20TO20(-219840), .W20TO21(-764147), .W20TO22(224877), .W20TO23(869767), .W20TO24(460398), .W20TO25(298423), .W20TO26(-779144), .W20TO27(161011), .W20TO28(-477341), .W20TO29(-212066), .W20TO30(-11421), .W20TO31(-390671), .W20TO32(953809), .W20TO33(-745992), .W20TO34(251836), .W20TO35(955421), .W20TO36(-157725), .W20TO37(37819), .W20TO38(-698411), .W20TO39(969544), .W20TO40(584802), .W20TO41(247307), .W20TO42(365680), .W20TO43(-933952), .W20TO44(281906), .W20TO45(358720), .W20TO46(719636), .W20TO47(287902), .W20TO48(8463), .W20TO49(777408), .W20TO50(531492), .W20TO51(-489842), .W20TO52(495045), .W20TO53(487524), .W20TO54(144972), .W20TO55(145529), .W20TO56(-173533), .W20TO57(810490), .W20TO58(739897), .W20TO59(360343), .W20TO60(868757), .W20TO61(658580), .W20TO62(81433), .W20TO63(-495238), .W21TO0(129517), .W21TO1(291665), .W21TO2(621452), .W21TO3(65567), .W21TO4(947670), .W21TO5(-583515), .W21TO6(-535366), .W21TO7(265650), .W21TO8(202589), .W21TO9(-377711), .W21TO10(273276), .W21TO11(943256), .W21TO12(829206), .W21TO13(601056), .W21TO14(-587670), .W21TO15(738225), .W21TO16(159392), .W21TO17(504588), .W21TO18(28080), .W21TO19(-833145), .W21TO20(-799539), .W21TO21(426780), .W21TO22(274560), .W21TO23(-510979), .W21TO24(-851833), .W21TO25(-744133), .W21TO26(552501), .W21TO27(-930545), .W21TO28(290353), .W21TO29(846169), .W21TO30(-782946), .W21TO31(884158), .W21TO32(357378), .W21TO33(-281636), .W21TO34(-615438), .W21TO35(226070), .W21TO36(13021), .W21TO37(-231526), .W21TO38(19795), .W21TO39(-7934), .W21TO40(865937), .W21TO41(-447383), .W21TO42(685496), .W21TO43(873465), .W21TO44(524169), .W21TO45(889514), .W21TO46(-660077), .W21TO47(-966283), .W21TO48(-10406), .W21TO49(-587301), .W21TO50(-393882), .W21TO51(531706), .W21TO52(-159974), .W21TO53(439320), .W21TO54(361116), .W21TO55(712032), .W21TO56(-231833), .W21TO57(876604), .W21TO58(921828), .W21TO59(23012), .W21TO60(-510363), .W21TO61(-620043), .W21TO62(17621), .W21TO63(-441478), .W22TO0(-782424), .W22TO1(-885973), .W22TO2(362797), .W22TO3(121597), .W22TO4(95144), .W22TO5(-733161), .W22TO6(687837), .W22TO7(-724225), .W22TO8(-372792), .W22TO9(473736), .W22TO10(-106921), .W22TO11(837745), .W22TO12(514015), .W22TO13(429359), .W22TO14(-544919), .W22TO15(-474090), .W22TO16(-298559), .W22TO17(838502), .W22TO18(311611), .W22TO19(700062), .W22TO20(-62779), .W22TO21(-778914), .W22TO22(-375683), .W22TO23(440260), .W22TO24(-656334), .W22TO25(-851123), .W22TO26(-993675), .W22TO27(-706532), .W22TO28(285250), .W22TO29(36350), .W22TO30(-212711), .W22TO31(-798715), .W22TO32(-574070), .W22TO33(810664), .W22TO34(-615973), .W22TO35(105344), .W22TO36(-203767), .W22TO37(-613625), .W22TO38(618742), .W22TO39(-613415), .W22TO40(862987), .W22TO41(-241258), .W22TO42(434948), .W22TO43(-824299), .W22TO44(-884460), .W22TO45(-587160), .W22TO46(-30526), .W22TO47(886095), .W22TO48(-711677), .W22TO49(990957), .W22TO50(-43574), .W22TO51(331027), .W22TO52(6829), .W22TO53(129681), .W22TO54(465527), .W22TO55(-459772), .W22TO56(563055), .W22TO57(-481346), .W22TO58(543109), .W22TO59(397356), .W22TO60(-21346), .W22TO61(848540), .W22TO62(-747618), .W22TO63(-976066), .W23TO0(693393), .W23TO1(-845307), .W23TO2(887070), .W23TO3(-847777), .W23TO4(-388870), .W23TO5(-639059), .W23TO6(-751979), .W23TO7(-594305), .W23TO8(436460), .W23TO9(310382), .W23TO10(25890), .W23TO11(-155234), .W23TO12(519570), .W23TO13(-24607), .W23TO14(831749), .W23TO15(544735), .W23TO16(423638), .W23TO17(-766809), .W23TO18(-313556), .W23TO19(-250112), .W23TO20(-74618), .W23TO21(-408242), .W23TO22(-434229), .W23TO23(938477), .W23TO24(-209817), .W23TO25(404895), .W23TO26(920049), .W23TO27(-181506), .W23TO28(327804), .W23TO29(683777), .W23TO30(-497247), .W23TO31(-579433), .W23TO32(-854080), .W23TO33(107500), .W23TO34(408083), .W23TO35(504672), .W23TO36(269618), .W23TO37(-874097), .W23TO38(-975641), .W23TO39(-553324), .W23TO40(-394952), .W23TO41(67441), .W23TO42(113848), .W23TO43(-357046), .W23TO44(330677), .W23TO45(-628564), .W23TO46(233148), .W23TO47(-291148), .W23TO48(-394531), .W23TO49(-518579), .W23TO50(331462), .W23TO51(-672568), .W23TO52(-861306), .W23TO53(-658591), .W23TO54(865341), .W23TO55(337825), .W23TO56(191598), .W23TO57(415966), .W23TO58(325437), .W23TO59(737115), .W23TO60(832309), .W23TO61(652981), .W23TO62(155380), .W23TO63(60525), .W24TO0(-707457), .W24TO1(204866), .W24TO2(-213955), .W24TO3(-903150), .W24TO4(519598), .W24TO5(333792), .W24TO6(-84627), .W24TO7(351159), .W24TO8(-149630), .W24TO9(535965), .W24TO10(851570), .W24TO11(-360937), .W24TO12(-407100), .W24TO13(-92638), .W24TO14(-566650), .W24TO15(-559190), .W24TO16(185230), .W24TO17(-404906), .W24TO18(-123519), .W24TO19(675605), .W24TO20(377856), .W24TO21(638200), .W24TO22(-590611), .W24TO23(715662), .W24TO24(83627), .W24TO25(853465), .W24TO26(-411434), .W24TO27(830988), .W24TO28(-842974), .W24TO29(-464871), .W24TO30(709221), .W24TO31(227784), .W24TO32(-39085), .W24TO33(376408), .W24TO34(-59297), .W24TO35(428403), .W24TO36(-103722), .W24TO37(-702150), .W24TO38(108691), .W24TO39(-220283), .W24TO40(248788), .W24TO41(961231), .W24TO42(-763025), .W24TO43(-63864), .W24TO44(-738272), .W24TO45(-63495), .W24TO46(-556334), .W24TO47(-214995), .W24TO48(759670), .W24TO49(-373520), .W24TO50(-572985), .W24TO51(757570), .W24TO52(-407673), .W24TO53(-748829), .W24TO54(-53400), .W24TO55(446940), .W24TO56(507328), .W24TO57(639938), .W24TO58(-996976), .W24TO59(-817152), .W24TO60(-984830), .W24TO61(498410), .W24TO62(719372), .W24TO63(-123240), .W25TO0(-945881), .W25TO1(828513), .W25TO2(-173589), .W25TO3(-169967), .W25TO4(386041), .W25TO5(874305), .W25TO6(231705), .W25TO7(383118), .W25TO8(470771), .W25TO9(-5549), .W25TO10(-280956), .W25TO11(-231752), .W25TO12(675984), .W25TO13(-793961), .W25TO14(664111), .W25TO15(-331346), .W25TO16(-286783), .W25TO17(-239580), .W25TO18(662201), .W25TO19(433828), .W25TO20(-806429), .W25TO21(-308769), .W25TO22(-926274), .W25TO23(564961), .W25TO24(-5432), .W25TO25(379385), .W25TO26(-847745), .W25TO27(819758), .W25TO28(268889), .W25TO29(780855), .W25TO30(-666242), .W25TO31(-329371), .W25TO32(-549875), .W25TO33(48874), .W25TO34(425286), .W25TO35(-310529), .W25TO36(748679), .W25TO37(-949467), .W25TO38(-413221), .W25TO39(4363), .W25TO40(377182), .W25TO41(-376866), .W25TO42(893498), .W25TO43(-511944), .W25TO44(-310219), .W25TO45(-311408), .W25TO46(-325853), .W25TO47(-885187), .W25TO48(-528278), .W25TO49(-149386), .W25TO50(-522604), .W25TO51(-423745), .W25TO52(564766), .W25TO53(322006), .W25TO54(52431), .W25TO55(319412), .W25TO56(837607), .W25TO57(741346), .W25TO58(853027), .W25TO59(-797772), .W25TO60(435638), .W25TO61(540145), .W25TO62(915205), .W25TO63(-947597), .W26TO0(-226371), .W26TO1(-536439), .W26TO2(-750876), .W26TO3(-818874), .W26TO4(69114), .W26TO5(723594), .W26TO6(-531775), .W26TO7(-174535), .W26TO8(-546999), .W26TO9(-123277), .W26TO10(390978), .W26TO11(396332), .W26TO12(411188), .W26TO13(-275071), .W26TO14(-882750), .W26TO15(243640), .W26TO16(-196205), .W26TO17(323677), .W26TO18(-468787), .W26TO19(913491), .W26TO20(-495600), .W26TO21(125010), .W26TO22(210565), .W26TO23(-144586), .W26TO24(632495), .W26TO25(101800), .W26TO26(29853), .W26TO27(-778112), .W26TO28(-448339), .W26TO29(598545), .W26TO30(714190), .W26TO31(-567446), .W26TO32(997090), .W26TO33(-903878), .W26TO34(-244136), .W26TO35(-864648), .W26TO36(-230075), .W26TO37(987134), .W26TO38(-810531), .W26TO39(-750454), .W26TO40(828933), .W26TO41(-293665), .W26TO42(-319596), .W26TO43(-146232), .W26TO44(327653), .W26TO45(144334), .W26TO46(-444248), .W26TO47(477984), .W26TO48(-395534), .W26TO49(721963), .W26TO50(233267), .W26TO51(-959031), .W26TO52(-462584), .W26TO53(-604243), .W26TO54(-281024), .W26TO55(283831), .W26TO56(-355396), .W26TO57(-856922), .W26TO58(835753), .W26TO59(-828328), .W26TO60(-828116), .W26TO61(666910), .W26TO62(-977215), .W26TO63(994260), .W27TO0(678598), .W27TO1(-405729), .W27TO2(-295675), .W27TO3(863532), .W27TO4(-753558), .W27TO5(106016), .W27TO6(585612), .W27TO7(-746782), .W27TO8(-108293), .W27TO9(-86638), .W27TO10(914182), .W27TO11(40831), .W27TO12(985442), .W27TO13(-885990), .W27TO14(-452259), .W27TO15(-430640), .W27TO16(464631), .W27TO17(-887553), .W27TO18(517966), .W27TO19(633102), .W27TO20(-65559), .W27TO21(-521662), .W27TO22(-387045), .W27TO23(410925), .W27TO24(-81252), .W27TO25(-551632), .W27TO26(444683), .W27TO27(607384), .W27TO28(824865), .W27TO29(199423), .W27TO30(479336), .W27TO31(-887218), .W27TO32(404152), .W27TO33(-278556), .W27TO34(-994037), .W27TO35(528021), .W27TO36(774541), .W27TO37(-513867), .W27TO38(-775709), .W27TO39(658532), .W27TO40(191431), .W27TO41(-448789), .W27TO42(831633), .W27TO43(-991321), .W27TO44(-157554), .W27TO45(-465691), .W27TO46(521224), .W27TO47(-745790), .W27TO48(461401), .W27TO49(-563660), .W27TO50(-996763), .W27TO51(426699), .W27TO52(-102468), .W27TO53(859878), .W27TO54(-668769), .W27TO55(146828), .W27TO56(199534), .W27TO57(-324164), .W27TO58(428617), .W27TO59(346153), .W27TO60(730031), .W27TO61(-933892), .W27TO62(267510), .W27TO63(584187), .W28TO0(934218), .W28TO1(-930596), .W28TO2(-207714), .W28TO3(339870), .W28TO4(696465), .W28TO5(-388600), .W28TO6(-362203), .W28TO7(569208), .W28TO8(-767404), .W28TO9(230880), .W28TO10(761494), .W28TO11(-102110), .W28TO12(74328), .W28TO13(130445), .W28TO14(-690734), .W28TO15(552161), .W28TO16(416832), .W28TO17(613912), .W28TO18(688321), .W28TO19(172455), .W28TO20(-692801), .W28TO21(415078), .W28TO22(-927072), .W28TO23(364841), .W28TO24(-497390), .W28TO25(-82347), .W28TO26(-273936), .W28TO27(-898336), .W28TO28(681033), .W28TO29(476842), .W28TO30(-203849), .W28TO31(564952), .W28TO32(80776), .W28TO33(865534), .W28TO34(668334), .W28TO35(-755546), .W28TO36(-34618), .W28TO37(-200141), .W28TO38(730641), .W28TO39(879915), .W28TO40(-547006), .W28TO41(-74869), .W28TO42(-814031), .W28TO43(390465), .W28TO44(627439), .W28TO45(-717997), .W28TO46(-703201), .W28TO47(206507), .W28TO48(869800), .W28TO49(-222990), .W28TO50(-428371), .W28TO51(-189035), .W28TO52(831182), .W28TO53(339923), .W28TO54(-406307), .W28TO55(208602), .W28TO56(357273), .W28TO57(-298160), .W28TO58(530388), .W28TO59(895417), .W28TO60(-631646), .W28TO61(-501615), .W28TO62(172071), .W28TO63(-435589), .W29TO0(792105), .W29TO1(522989), .W29TO2(-448235), .W29TO3(875158), .W29TO4(291874), .W29TO5(634394), .W29TO6(-53840), .W29TO7(596836), .W29TO8(-369071), .W29TO9(465636), .W29TO10(-11687), .W29TO11(-648356), .W29TO12(-958169), .W29TO13(-964649), .W29TO14(868087), .W29TO15(204357), .W29TO16(578913), .W29TO17(518176), .W29TO18(-688155), .W29TO19(-12834), .W29TO20(684306), .W29TO21(-879072), .W29TO22(-793455), .W29TO23(329446), .W29TO24(743549), .W29TO25(-842651), .W29TO26(722159), .W29TO27(198503), .W29TO28(751751), .W29TO29(-405010), .W29TO30(-390820), .W29TO31(924932), .W29TO32(-395211), .W29TO33(-310855), .W29TO34(-435642), .W29TO35(-896309), .W29TO36(468453), .W29TO37(-136187), .W29TO38(546373), .W29TO39(473988), .W29TO40(462057), .W29TO41(604148), .W29TO42(-733959), .W29TO43(28432), .W29TO44(279673), .W29TO45(786510), .W29TO46(610664), .W29TO47(-435952), .W29TO48(-553889), .W29TO49(806410), .W29TO50(-401575), .W29TO51(-493990), .W29TO52(-888598), .W29TO53(993007), .W29TO54(618078), .W29TO55(567507), .W29TO56(-938139), .W29TO57(62687), .W29TO58(66585), .W29TO59(566158), .W29TO60(689209), .W29TO61(704075), .W29TO62(-54585), .W29TO63(589771), .W30TO0(948863), .W30TO1(-879067), .W30TO2(739202), .W30TO3(-262806), .W30TO4(-140320), .W30TO5(-984263), .W30TO6(309986), .W30TO7(172559), .W30TO8(979592), .W30TO9(477543), .W30TO10(27541), .W30TO11(143), .W30TO12(502260), .W30TO13(-811574), .W30TO14(928407), .W30TO15(-663941), .W30TO16(-408250), .W30TO17(-744603), .W30TO18(111912), .W30TO19(-632615), .W30TO20(-516114), .W30TO21(-963901), .W30TO22(-665276), .W30TO23(-164469), .W30TO24(21880), .W30TO25(-506069), .W30TO26(238762), .W30TO27(-397422), .W30TO28(473542), .W30TO29(-70187), .W30TO30(739038), .W30TO31(604314), .W30TO32(-472596), .W30TO33(330949), .W30TO34(-231676), .W30TO35(-405644), .W30TO36(596966), .W30TO37(400364), .W30TO38(-794687), .W30TO39(-947932), .W30TO40(-534971), .W30TO41(938390), .W30TO42(527989), .W30TO43(551318), .W30TO44(-963507), .W30TO45(-541485), .W30TO46(-594020), .W30TO47(690833), .W30TO48(858787), .W30TO49(-814896), .W30TO50(-18231), .W30TO51(490601), .W30TO52(457611), .W30TO53(346129), .W30TO54(-226615), .W30TO55(432224), .W30TO56(763813), .W30TO57(65438), .W30TO58(-427940), .W30TO59(724383), .W30TO60(789030), .W30TO61(-329914), .W30TO62(979380), .W30TO63(188088), .W31TO0(837270), .W31TO1(-152721), .W31TO2(243322), .W31TO3(-396142), .W31TO4(178238), .W31TO5(-591882), .W31TO6(-592748), .W31TO7(424849), .W31TO8(-35817), .W31TO9(-132114), .W31TO10(-611827), .W31TO11(929765), .W31TO12(473699), .W31TO13(-450170), .W31TO14(-61834), .W31TO15(-638309), .W31TO16(799296), .W31TO17(482352), .W31TO18(326690), .W31TO19(-948424), .W31TO20(-59061), .W31TO21(-926782), .W31TO22(-993986), .W31TO23(633491), .W31TO24(-554160), .W31TO25(-230845), .W31TO26(-820455), .W31TO27(64604), .W31TO28(759716), .W31TO29(-163109), .W31TO30(761698), .W31TO31(-82321), .W31TO32(905151), .W31TO33(-391131), .W31TO34(-740325), .W31TO35(97535), .W31TO36(-534207), .W31TO37(-488562), .W31TO38(2921), .W31TO39(-922952), .W31TO40(-602243), .W31TO41(-71438), .W31TO42(460841), .W31TO43(-223512), .W31TO44(470373), .W31TO45(-994221), .W31TO46(-192370), .W31TO47(-512295), .W31TO48(-926305), .W31TO49(-895516), .W31TO50(-255003), .W31TO51(-143108), .W31TO52(284686), .W31TO53(658620), .W31TO54(-688295), .W31TO55(496573), .W31TO56(-562408), .W31TO57(-782197), .W31TO58(894259), .W31TO59(475605), .W31TO60(57850), .W31TO61(610874), .W31TO62(309474), .W31TO63(87499), .W32TO0(-428722), .W32TO1(-139354), .W32TO2(589363), .W32TO3(-943812), .W32TO4(442825), .W32TO5(422861), .W32TO6(169322), .W32TO7(489545), .W32TO8(297326), .W32TO9(687712), .W32TO10(-297515), .W32TO11(332300), .W32TO12(419207), .W32TO13(-744265), .W32TO14(-748348), .W32TO15(840266), .W32TO16(-573743), .W32TO17(-357166), .W32TO18(-692402), .W32TO19(-324545), .W32TO20(568248), .W32TO21(400147), .W32TO22(422376), .W32TO23(696173), .W32TO24(974336), .W32TO25(-273108), .W32TO26(-388174), .W32TO27(-168000), .W32TO28(-27102), .W32TO29(968858), .W32TO30(529401), .W32TO31(162483), .W32TO32(-720232), .W32TO33(816414), .W32TO34(-575656), .W32TO35(857112), .W32TO36(-357712), .W32TO37(-364289), .W32TO38(-28560), .W32TO39(-525046), .W32TO40(727921), .W32TO41(766967), .W32TO42(652609), .W32TO43(-447749), .W32TO44(82325), .W32TO45(739893), .W32TO46(-598969), .W32TO47(-497238), .W32TO48(-876015), .W32TO49(-823373), .W32TO50(-386248), .W32TO51(-154312), .W32TO52(672862), .W32TO53(394768), .W32TO54(866538), .W32TO55(530568), .W32TO56(341136), .W32TO57(-589804), .W32TO58(-518051), .W32TO59(109553), .W32TO60(611663), .W32TO61(-547944), .W32TO62(-461156), .W32TO63(330683), .W33TO0(158063), .W33TO1(418219), .W33TO2(686544), .W33TO3(-753292), .W33TO4(-543974), .W33TO5(-286182), .W33TO6(-787592), .W33TO7(-483784), .W33TO8(-790991), .W33TO9(-536875), .W33TO10(466793), .W33TO11(-329709), .W33TO12(28356), .W33TO13(367871), .W33TO14(665633), .W33TO15(-852493), .W33TO16(251105), .W33TO17(-626179), .W33TO18(823749), .W33TO19(-188925), .W33TO20(-21454), .W33TO21(-111305), .W33TO22(650329), .W33TO23(533193), .W33TO24(200125), .W33TO25(769869), .W33TO26(-546785), .W33TO27(175608), .W33TO28(86748), .W33TO29(-859625), .W33TO30(69906), .W33TO31(-897547), .W33TO32(-151876), .W33TO33(-556714), .W33TO34(524361), .W33TO35(58645), .W33TO36(-96812), .W33TO37(138411), .W33TO38(-848877), .W33TO39(506563), .W33TO40(732661), .W33TO41(495453), .W33TO42(256350), .W33TO43(-991928), .W33TO44(-826385), .W33TO45(-957900), .W33TO46(193295), .W33TO47(92972), .W33TO48(-498021), .W33TO49(582583), .W33TO50(-662985), .W33TO51(-193118), .W33TO52(-210818), .W33TO53(736684), .W33TO54(-999798), .W33TO55(164291), .W33TO56(348737), .W33TO57(361788), .W33TO58(-869922), .W33TO59(-708555), .W33TO60(155232), .W33TO61(427985), .W33TO62(-575904), .W33TO63(660468), .W34TO0(-626395), .W34TO1(-535080), .W34TO2(-840612), .W34TO3(-632742), .W34TO4(-168043), .W34TO5(-672338), .W34TO6(140132), .W34TO7(486410), .W34TO8(-369092), .W34TO9(-11415), .W34TO10(-197527), .W34TO11(-744498), .W34TO12(-819022), .W34TO13(771289), .W34TO14(-926553), .W34TO15(23190), .W34TO16(-461276), .W34TO17(773441), .W34TO18(-248764), .W34TO19(-595442), .W34TO20(651800), .W34TO21(-140154), .W34TO22(-534299), .W34TO23(183935), .W34TO24(-634202), .W34TO25(787079), .W34TO26(116762), .W34TO27(-99779), .W34TO28(-618060), .W34TO29(-662951), .W34TO30(-405807), .W34TO31(-375076), .W34TO32(25527), .W34TO33(-540780), .W34TO34(169457), .W34TO35(735418), .W34TO36(-709011), .W34TO37(529683), .W34TO38(207568), .W34TO39(-294459), .W34TO40(157061), .W34TO41(645001), .W34TO42(-891838), .W34TO43(418922), .W34TO44(789865), .W34TO45(-500134), .W34TO46(-385548), .W34TO47(-881755), .W34TO48(-746155), .W34TO49(200556), .W34TO50(855140), .W34TO51(-678664), .W34TO52(479956), .W34TO53(83827), .W34TO54(-468691), .W34TO55(-141158), .W34TO56(78525), .W34TO57(374672), .W34TO58(-489060), .W34TO59(-48875), .W34TO60(780930), .W34TO61(-657052), .W34TO62(-143332), .W34TO63(486546), .W35TO0(521403), .W35TO1(-204250), .W35TO2(-233920), .W35TO3(-43858), .W35TO4(-437591), .W35TO5(177627), .W35TO6(248746), .W35TO7(-99999), .W35TO8(-112840), .W35TO9(-789701), .W35TO10(698401), .W35TO11(257674), .W35TO12(-581693), .W35TO13(909858), .W35TO14(314943), .W35TO15(179554), .W35TO16(125923), .W35TO17(795614), .W35TO18(929551), .W35TO19(-507799), .W35TO20(350415), .W35TO21(-816926), .W35TO22(138293), .W35TO23(527606), .W35TO24(-545356), .W35TO25(493271), .W35TO26(996882), .W35TO27(-377454), .W35TO28(-81176), .W35TO29(952473), .W35TO30(687899), .W35TO31(557539), .W35TO32(326588), .W35TO33(-595225), .W35TO34(249843), .W35TO35(409), .W35TO36(-488233), .W35TO37(-395650), .W35TO38(-192286), .W35TO39(-848304), .W35TO40(-932855), .W35TO41(753562), .W35TO42(371248), .W35TO43(-494544), .W35TO44(-485447), .W35TO45(207712), .W35TO46(-352610), .W35TO47(91174), .W35TO48(-517913), .W35TO49(726788), .W35TO50(778084), .W35TO51(406380), .W35TO52(-82803), .W35TO53(457879), .W35TO54(-545905), .W35TO55(523312), .W35TO56(499666), .W35TO57(77668), .W35TO58(885285), .W35TO59(137375), .W35TO60(-48475), .W35TO61(494908), .W35TO62(673916), .W35TO63(-299971), .W36TO0(67894), .W36TO1(-434884), .W36TO2(-574405), .W36TO3(539506), .W36TO4(-245536), .W36TO5(-535059), .W36TO6(968843), .W36TO7(-120145), .W36TO8(-883513), .W36TO9(424253), .W36TO10(-844131), .W36TO11(133773), .W36TO12(296904), .W36TO13(148891), .W36TO14(58930), .W36TO15(4371), .W36TO16(-584568), .W36TO17(301249), .W36TO18(-698716), .W36TO19(-763186), .W36TO20(-685908), .W36TO21(395464), .W36TO22(-578722), .W36TO23(-35652), .W36TO24(-854329), .W36TO25(922468), .W36TO26(-468823), .W36TO27(646865), .W36TO28(754259), .W36TO29(-275456), .W36TO30(665450), .W36TO31(-219989), .W36TO32(-622584), .W36TO33(663638), .W36TO34(-462479), .W36TO35(261410), .W36TO36(197692), .W36TO37(726256), .W36TO38(-816795), .W36TO39(-344571), .W36TO40(364913), .W36TO41(-260516), .W36TO42(136335), .W36TO43(-854634), .W36TO44(-88937), .W36TO45(-829928), .W36TO46(884304), .W36TO47(628109), .W36TO48(-819303), .W36TO49(93199), .W36TO50(-996444), .W36TO51(572117), .W36TO52(275445), .W36TO53(677956), .W36TO54(-608984), .W36TO55(-203706), .W36TO56(440639), .W36TO57(389894), .W36TO58(-17265), .W36TO59(-428573), .W36TO60(349393), .W36TO61(977869), .W36TO62(-861403), .W36TO63(92972), .W37TO0(11393), .W37TO1(455874), .W37TO2(866136), .W37TO3(-480294), .W37TO4(-388517), .W37TO5(469933), .W37TO6(881567), .W37TO7(216548), .W37TO8(705726), .W37TO9(-534310), .W37TO10(450391), .W37TO11(251268), .W37TO12(349662), .W37TO13(-809667), .W37TO14(808964), .W37TO15(165383), .W37TO16(-341503), .W37TO17(308104), .W37TO18(-305443), .W37TO19(-697345), .W37TO20(-481755), .W37TO21(-16558), .W37TO22(474606), .W37TO23(-508076), .W37TO24(44614), .W37TO25(894183), .W37TO26(-871084), .W37TO27(-949001), .W37TO28(-236526), .W37TO29(-600241), .W37TO30(285814), .W37TO31(-543013), .W37TO32(239284), .W37TO33(738900), .W37TO34(-779165), .W37TO35(22373), .W37TO36(-942016), .W37TO37(414936), .W37TO38(-673826), .W37TO39(261022), .W37TO40(-924942), .W37TO41(902036), .W37TO42(-134928), .W37TO43(-769737), .W37TO44(352764), .W37TO45(774649), .W37TO46(-464144), .W37TO47(-154134), .W37TO48(727684), .W37TO49(494954), .W37TO50(-191964), .W37TO51(-327247), .W37TO52(-839592), .W37TO53(56125), .W37TO54(-958977), .W37TO55(-374751), .W37TO56(42642), .W37TO57(398430), .W37TO58(-833362), .W37TO59(240913), .W37TO60(-685257), .W37TO61(930356), .W37TO62(-742388), .W37TO63(8664), .W38TO0(-937206), .W38TO1(-24398), .W38TO2(-113882), .W38TO3(-671605), .W38TO4(-345453), .W38TO5(817517), .W38TO6(545241), .W38TO7(-230595), .W38TO8(-759460), .W38TO9(-372700), .W38TO10(-588373), .W38TO11(-95116), .W38TO12(-964054), .W38TO13(-937342), .W38TO14(-246320), .W38TO15(245131), .W38TO16(160797), .W38TO17(-459313), .W38TO18(593765), .W38TO19(-251407), .W38TO20(-234334), .W38TO21(542115), .W38TO22(-238857), .W38TO23(663163), .W38TO24(968002), .W38TO25(-29537), .W38TO26(7834), .W38TO27(638570), .W38TO28(-402983), .W38TO29(-553252), .W38TO30(-159445), .W38TO31(589706), .W38TO32(104137), .W38TO33(670491), .W38TO34(498980), .W38TO35(511944), .W38TO36(-100145), .W38TO37(-485960), .W38TO38(658818), .W38TO39(843721), .W38TO40(-897112), .W38TO41(142612), .W38TO42(-809062), .W38TO43(390366), .W38TO44(-756237), .W38TO45(875937), .W38TO46(-37835), .W38TO47(475687), .W38TO48(681363), .W38TO49(-557902), .W38TO50(-78668), .W38TO51(-307883), .W38TO52(-345054), .W38TO53(614134), .W38TO54(-654273), .W38TO55(603354), .W38TO56(-121533), .W38TO57(186903), .W38TO58(659080), .W38TO59(746998), .W38TO60(-844836), .W38TO61(-969980), .W38TO62(-986518), .W38TO63(344737), .W39TO0(-902110), .W39TO1(713734), .W39TO2(-229315), .W39TO3(-246433), .W39TO4(767768), .W39TO5(419147), .W39TO6(55187), .W39TO7(-869972), .W39TO8(80706), .W39TO9(503310), .W39TO10(421330), .W39TO11(-925476), .W39TO12(768456), .W39TO13(317794), .W39TO14(435697), .W39TO15(610590), .W39TO16(-345409), .W39TO17(295425), .W39TO18(-202579), .W39TO19(-64871), .W39TO20(451741), .W39TO21(858670), .W39TO22(-289778), .W39TO23(394352), .W39TO24(953933), .W39TO25(805289), .W39TO26(938762), .W39TO27(-803224), .W39TO28(-658747), .W39TO29(432344), .W39TO30(-20111), .W39TO31(430098), .W39TO32(463905), .W39TO33(768643), .W39TO34(-474336), .W39TO35(-913515), .W39TO36(-923735), .W39TO37(812871), .W39TO38(139063), .W39TO39(868566), .W39TO40(754677), .W39TO41(541670), .W39TO42(437752), .W39TO43(-947397), .W39TO44(-993954), .W39TO45(972346), .W39TO46(-567538), .W39TO47(-748213), .W39TO48(-55167), .W39TO49(-293161), .W39TO50(-691357), .W39TO51(856822), .W39TO52(46277), .W39TO53(-44246), .W39TO54(-742255), .W39TO55(-673738), .W39TO56(-197763), .W39TO57(405559), .W39TO58(-649107), .W39TO59(861996), .W39TO60(755675), .W39TO61(-385815), .W39TO62(490368), .W39TO63(837574), .W40TO0(-102617), .W40TO1(-111875), .W40TO2(-628935), .W40TO3(-688582), .W40TO4(-332218), .W40TO5(-27139), .W40TO6(-769722), .W40TO7(92936), .W40TO8(-450293), .W40TO9(684453), .W40TO10(273925), .W40TO11(-145077), .W40TO12(38205), .W40TO13(675462), .W40TO14(-182605), .W40TO15(-637227), .W40TO16(599876), .W40TO17(-686020), .W40TO18(650669), .W40TO19(-823040), .W40TO20(-314069), .W40TO21(135612), .W40TO22(726348), .W40TO23(305481), .W40TO24(-744340), .W40TO25(726126), .W40TO26(-770688), .W40TO27(-757549), .W40TO28(988715), .W40TO29(-656647), .W40TO30(-272401), .W40TO31(138302), .W40TO32(513201), .W40TO33(-667017), .W40TO34(836877), .W40TO35(-14882), .W40TO36(-606909), .W40TO37(-64827), .W40TO38(-707033), .W40TO39(-651612), .W40TO40(450197), .W40TO41(-813832), .W40TO42(-682089), .W40TO43(-658958), .W40TO44(346347), .W40TO45(750183), .W40TO46(9270), .W40TO47(-495774), .W40TO48(226939), .W40TO49(752090), .W40TO50(-944283), .W40TO51(-547927), .W40TO52(271077), .W40TO53(619872), .W40TO54(129393), .W40TO55(-620070), .W40TO56(207641), .W40TO57(535027), .W40TO58(-491610), .W40TO59(-11181), .W40TO60(199278), .W40TO61(562289), .W40TO62(434413), .W40TO63(-257174), .W41TO0(-688861), .W41TO1(-143055), .W41TO2(-564348), .W41TO3(-669399), .W41TO4(-648722), .W41TO5(-516509), .W41TO6(754612), .W41TO7(116252), .W41TO8(-315930), .W41TO9(-335226), .W41TO10(160401), .W41TO11(-784769), .W41TO12(606206), .W41TO13(628472), .W41TO14(800411), .W41TO15(416397), .W41TO16(106298), .W41TO17(907560), .W41TO18(259634), .W41TO19(-865991), .W41TO20(817156), .W41TO21(504921), .W41TO22(-595846), .W41TO23(77507), .W41TO24(952480), .W41TO25(187255), .W41TO26(873375), .W41TO27(-506974), .W41TO28(405155), .W41TO29(-847416), .W41TO30(583053), .W41TO31(-966152), .W41TO32(-135331), .W41TO33(763215), .W41TO34(-191935), .W41TO35(891076), .W41TO36(183198), .W41TO37(-231918), .W41TO38(503045), .W41TO39(-796772), .W41TO40(-467858), .W41TO41(-890600), .W41TO42(109279), .W41TO43(122253), .W41TO44(814444), .W41TO45(84690), .W41TO46(389162), .W41TO47(-377695), .W41TO48(-58950), .W41TO49(-308544), .W41TO50(-596167), .W41TO51(-544939), .W41TO52(-572097), .W41TO53(865467), .W41TO54(993558), .W41TO55(-40658), .W41TO56(580610), .W41TO57(-119751), .W41TO58(-497091), .W41TO59(-896586), .W41TO60(954317), .W41TO61(366284), .W41TO62(-28763), .W41TO63(691294), .W42TO0(414903), .W42TO1(274330), .W42TO2(-296347), .W42TO3(-171342), .W42TO4(403471), .W42TO5(32846), .W42TO6(-844673), .W42TO7(575672), .W42TO8(651423), .W42TO9(546492), .W42TO10(650174), .W42TO11(-253972), .W42TO12(198469), .W42TO13(-469452), .W42TO14(-645484), .W42TO15(-515218), .W42TO16(754127), .W42TO17(-617093), .W42TO18(507222), .W42TO19(125515), .W42TO20(876335), .W42TO21(926643), .W42TO22(910978), .W42TO23(-599028), .W42TO24(787049), .W42TO25(-857654), .W42TO26(-328108), .W42TO27(-907748), .W42TO28(-69185), .W42TO29(447054), .W42TO30(983900), .W42TO31(-395345), .W42TO32(-710019), .W42TO33(616499), .W42TO34(-798904), .W42TO35(172560), .W42TO36(-871302), .W42TO37(-274223), .W42TO38(406886), .W42TO39(-775006), .W42TO40(191574), .W42TO41(-611957), .W42TO42(534665), .W42TO43(783681), .W42TO44(393067), .W42TO45(518014), .W42TO46(-200171), .W42TO47(-353792), .W42TO48(41303), .W42TO49(295184), .W42TO50(-611457), .W42TO51(-353808), .W42TO52(353972), .W42TO53(-901256), .W42TO54(-884489), .W42TO55(350505), .W42TO56(690393), .W42TO57(341723), .W42TO58(18088), .W42TO59(-524661), .W42TO60(-673176), .W42TO61(-690711), .W42TO62(-493518), .W42TO63(71285), .W43TO0(962770), .W43TO1(-694148), .W43TO2(187095), .W43TO3(475391), .W43TO4(808389), .W43TO5(-799810), .W43TO6(-26646), .W43TO7(246477), .W43TO8(844549), .W43TO9(-424565), .W43TO10(-139377), .W43TO11(-989736), .W43TO12(217089), .W43TO13(396421), .W43TO14(-494516), .W43TO15(917631), .W43TO16(187390), .W43TO17(-928384), .W43TO18(-29114), .W43TO19(282893), .W43TO20(-176866), .W43TO21(-58776), .W43TO22(899203), .W43TO23(-651672), .W43TO24(467809), .W43TO25(-40379), .W43TO26(435528), .W43TO27(-32546), .W43TO28(-448821), .W43TO29(-601687), .W43TO30(791232), .W43TO31(832217), .W43TO32(430839), .W43TO33(198845), .W43TO34(-618620), .W43TO35(75032), .W43TO36(-851334), .W43TO37(-343614), .W43TO38(533055), .W43TO39(356283), .W43TO40(-800965), .W43TO41(-618934), .W43TO42(-583825), .W43TO43(724640), .W43TO44(787574), .W43TO45(-570704), .W43TO46(-257527), .W43TO47(238754), .W43TO48(-345584), .W43TO49(747209), .W43TO50(-661252), .W43TO51(369097), .W43TO52(-727850), .W43TO53(-531661), .W43TO54(45694), .W43TO55(771775), .W43TO56(637745), .W43TO57(-430378), .W43TO58(356173), .W43TO59(-774338), .W43TO60(-68802), .W43TO61(566254), .W43TO62(771037), .W43TO63(948658), .W44TO0(692475), .W44TO1(243082), .W44TO2(677177), .W44TO3(-502909), .W44TO4(222908), .W44TO5(-104842), .W44TO6(-681912), .W44TO7(-223212), .W44TO8(-735062), .W44TO9(824341), .W44TO10(-378443), .W44TO11(-942925), .W44TO12(-339619), .W44TO13(-526441), .W44TO14(-423433), .W44TO15(-872719), .W44TO16(-838160), .W44TO17(290211), .W44TO18(212863), .W44TO19(269855), .W44TO20(-308061), .W44TO21(31500), .W44TO22(470590), .W44TO23(241234), .W44TO24(358107), .W44TO25(943966), .W44TO26(-467900), .W44TO27(-820341), .W44TO28(131902), .W44TO29(700227), .W44TO30(941926), .W44TO31(-153724), .W44TO32(-659030), .W44TO33(-641809), .W44TO34(-935437), .W44TO35(-800005), .W44TO36(591548), .W44TO37(-580921), .W44TO38(-215986), .W44TO39(-952746), .W44TO40(-874531), .W44TO41(190650), .W44TO42(-251139), .W44TO43(-238710), .W44TO44(598575), .W44TO45(-363534), .W44TO46(260868), .W44TO47(679069), .W44TO48(-33601), .W44TO49(-292052), .W44TO50(-125502), .W44TO51(773607), .W44TO52(741094), .W44TO53(-356523), .W44TO54(452355), .W44TO55(-37035), .W44TO56(63313), .W44TO57(461166), .W44TO58(485336), .W44TO59(-106089), .W44TO60(195158), .W44TO61(-508223), .W44TO62(195272), .W44TO63(-222719), .W45TO0(-905839), .W45TO1(563387), .W45TO2(-877346), .W45TO3(117021), .W45TO4(-217206), .W45TO5(-916340), .W45TO6(-884883), .W45TO7(-836858), .W45TO8(625257), .W45TO9(-5651), .W45TO10(6808), .W45TO11(-938410), .W45TO12(964785), .W45TO13(-846635), .W45TO14(959966), .W45TO15(138393), .W45TO16(-895278), .W45TO17(923643), .W45TO18(826198), .W45TO19(976465), .W45TO20(831525), .W45TO21(963490), .W45TO22(-752048), .W45TO23(-627114), .W45TO24(169376), .W45TO25(-862910), .W45TO26(639402), .W45TO27(-548187), .W45TO28(-241708), .W45TO29(-114634), .W45TO30(519566), .W45TO31(308853), .W45TO32(41775), .W45TO33(892129), .W45TO34(107525), .W45TO35(530318), .W45TO36(-114189), .W45TO37(-300448), .W45TO38(-794302), .W45TO39(-789769), .W45TO40(81263), .W45TO41(-504708), .W45TO42(-969004), .W45TO43(-633375), .W45TO44(276616), .W45TO45(-807176), .W45TO46(601345), .W45TO47(-979660), .W45TO48(-498601), .W45TO49(445022), .W45TO50(-789627), .W45TO51(803557), .W45TO52(443631), .W45TO53(769407), .W45TO54(-618971), .W45TO55(-28790), .W45TO56(778632), .W45TO57(-446689), .W45TO58(-518452), .W45TO59(57838), .W45TO60(778283), .W45TO61(982022), .W45TO62(-204157), .W45TO63(-402082), .W46TO0(156046), .W46TO1(793583), .W46TO2(-603820), .W46TO3(822959), .W46TO4(-779480), .W46TO5(687524), .W46TO6(-817354), .W46TO7(-637238), .W46TO8(839419), .W46TO9(565864), .W46TO10(-959441), .W46TO11(477081), .W46TO12(-910608), .W46TO13(-97248), .W46TO14(413786), .W46TO15(-97598), .W46TO16(956935), .W46TO17(-753978), .W46TO18(-549984), .W46TO19(-750244), .W46TO20(-610172), .W46TO21(-765251), .W46TO22(-353771), .W46TO23(964481), .W46TO24(-887540), .W46TO25(50399), .W46TO26(652727), .W46TO27(923376), .W46TO28(267942), .W46TO29(632297), .W46TO30(950081), .W46TO31(626113), .W46TO32(233692), .W46TO33(2854), .W46TO34(-574130), .W46TO35(-673445), .W46TO36(-71050), .W46TO37(733035), .W46TO38(-941657), .W46TO39(870999), .W46TO40(740280), .W46TO41(-535657), .W46TO42(679263), .W46TO43(-23216), .W46TO44(543450), .W46TO45(357684), .W46TO46(-195495), .W46TO47(144067), .W46TO48(70805), .W46TO49(724294), .W46TO50(255526), .W46TO51(125518), .W46TO52(885154), .W46TO53(-979456), .W46TO54(526166), .W46TO55(564136), .W46TO56(-806264), .W46TO57(470231), .W46TO58(698675), .W46TO59(712772), .W46TO60(-442268), .W46TO61(449954), .W46TO62(-525473), .W46TO63(-973328), .W47TO0(849318), .W47TO1(-132952), .W47TO2(382288), .W47TO3(190399), .W47TO4(-360785), .W47TO5(968684), .W47TO6(-935293), .W47TO7(473356), .W47TO8(-888379), .W47TO9(-573348), .W47TO10(-169972), .W47TO11(-70786), .W47TO12(630580), .W47TO13(-918904), .W47TO14(-980457), .W47TO15(-446191), .W47TO16(125499), .W47TO17(946569), .W47TO18(866370), .W47TO19(-59612), .W47TO20(-910510), .W47TO21(-135288), .W47TO22(595169), .W47TO23(699437), .W47TO24(-321574), .W47TO25(411397), .W47TO26(971360), .W47TO27(870538), .W47TO28(-300096), .W47TO29(765119), .W47TO30(432840), .W47TO31(741445), .W47TO32(-35704), .W47TO33(983909), .W47TO34(-553686), .W47TO35(-506623), .W47TO36(854212), .W47TO37(863784), .W47TO38(-540582), .W47TO39(696687), .W47TO40(209509), .W47TO41(-625387), .W47TO42(99295), .W47TO43(640522), .W47TO44(-254271), .W47TO45(220493), .W47TO46(-462414), .W47TO47(-754273), .W47TO48(502793), .W47TO49(-953904), .W47TO50(-214871), .W47TO51(-468058), .W47TO52(817786), .W47TO53(-394539), .W47TO54(71339), .W47TO55(-484372), .W47TO56(341420), .W47TO57(803462), .W47TO58(92492), .W47TO59(442087), .W47TO60(464775), .W47TO61(-418970), .W47TO62(-394224), .W47TO63(774558), .W48TO0(-893489), .W48TO1(-471665), .W48TO2(-78701), .W48TO3(-567128), .W48TO4(274705), .W48TO5(843312), .W48TO6(764884), .W48TO7(253505), .W48TO8(843817), .W48TO9(162943), .W48TO10(489789), .W48TO11(287146), .W48TO12(20852), .W48TO13(450504), .W48TO14(-614396), .W48TO15(724145), .W48TO16(-637654), .W48TO17(-355498), .W48TO18(-126309), .W48TO19(-342842), .W48TO20(-81745), .W48TO21(-327282), .W48TO22(766205), .W48TO23(-429096), .W48TO24(249156), .W48TO25(-702160), .W48TO26(-362936), .W48TO27(820184), .W48TO28(-196032), .W48TO29(-612348), .W48TO30(-839852), .W48TO31(13788), .W48TO32(-40748), .W48TO33(584347), .W48TO34(-437561), .W48TO35(300608), .W48TO36(40175), .W48TO37(-537636), .W48TO38(-728268), .W48TO39(-610329), .W48TO40(602217), .W48TO41(245951), .W48TO42(-943145), .W48TO43(592695), .W48TO44(-474810), .W48TO45(433431), .W48TO46(663790), .W48TO47(-962789), .W48TO48(-74200), .W48TO49(-385996), .W48TO50(669417), .W48TO51(-737854), .W48TO52(855418), .W48TO53(-939523), .W48TO54(679081), .W48TO55(557504), .W48TO56(-143558), .W48TO57(-746176), .W48TO58(-196958), .W48TO59(471936), .W48TO60(-492216), .W48TO61(973314), .W48TO62(-339818), .W48TO63(-907462), .W49TO0(52027), .W49TO1(7523), .W49TO2(-146125), .W49TO3(-388694), .W49TO4(944188), .W49TO5(331456), .W49TO6(43944), .W49TO7(659831), .W49TO8(365745), .W49TO9(-317602), .W49TO10(-210121), .W49TO11(231289), .W49TO12(874962), .W49TO13(-25638), .W49TO14(-157401), .W49TO15(-303425), .W49TO16(-770705), .W49TO17(-786380), .W49TO18(-990254), .W49TO19(531552), .W49TO20(-324420), .W49TO21(-214095), .W49TO22(-685558), .W49TO23(709524), .W49TO24(832159), .W49TO25(-780219), .W49TO26(-880225), .W49TO27(343678), .W49TO28(688471), .W49TO29(808701), .W49TO30(240411), .W49TO31(-733977), .W49TO32(714778), .W49TO33(-637106), .W49TO34(-406688), .W49TO35(719783), .W49TO36(527671), .W49TO37(820225), .W49TO38(-861658), .W49TO39(278080), .W49TO40(-381904), .W49TO41(993343), .W49TO42(-247639), .W49TO43(-682233), .W49TO44(-102846), .W49TO45(-24595), .W49TO46(-706498), .W49TO47(-457240), .W49TO48(157211), .W49TO49(950734), .W49TO50(815544), .W49TO51(453810), .W49TO52(-625871), .W49TO53(352373), .W49TO54(-648889), .W49TO55(15056), .W49TO56(-672441), .W49TO57(664180), .W49TO58(970723), .W49TO59(-994248), .W49TO60(-114556), .W49TO61(-852701), .W49TO62(-146595), .W49TO63(-831019), .W50TO0(-523287), .W50TO1(720332), .W50TO2(441986), .W50TO3(-272408), .W50TO4(-782012), .W50TO5(74750), .W50TO6(608115), .W50TO7(345947), .W50TO8(-25707), .W50TO9(-679317), .W50TO10(-963724), .W50TO11(-557043), .W50TO12(707849), .W50TO13(-496503), .W50TO14(-518462), .W50TO15(506329), .W50TO16(157266), .W50TO17(-747012), .W50TO18(379999), .W50TO19(949296), .W50TO20(800675), .W50TO21(-758991), .W50TO22(342335), .W50TO23(-63595), .W50TO24(120867), .W50TO25(116005), .W50TO26(-818560), .W50TO27(-508282), .W50TO28(557616), .W50TO29(27849), .W50TO30(174151), .W50TO31(974238), .W50TO32(376900), .W50TO33(-956637), .W50TO34(416834), .W50TO35(-68413), .W50TO36(-59752), .W50TO37(-490027), .W50TO38(544547), .W50TO39(-409003), .W50TO40(-320950), .W50TO41(-82476), .W50TO42(-23074), .W50TO43(429676), .W50TO44(-793629), .W50TO45(-477967), .W50TO46(332343), .W50TO47(298067), .W50TO48(-21702), .W50TO49(459149), .W50TO50(60082), .W50TO51(180877), .W50TO52(-390760), .W50TO53(106139), .W50TO54(10839), .W50TO55(-997918), .W50TO56(-557210), .W50TO57(-294596), .W50TO58(-156031), .W50TO59(-642243), .W50TO60(-488212), .W50TO61(713155), .W50TO62(615195), .W50TO63(449884), .W51TO0(-848978), .W51TO1(759465), .W51TO2(706123), .W51TO3(-598404), .W51TO4(-502386), .W51TO5(860213), .W51TO6(403103), .W51TO7(63916), .W51TO8(-493822), .W51TO9(134102), .W51TO10(-190178), .W51TO11(-371555), .W51TO12(-384973), .W51TO13(-306784), .W51TO14(74360), .W51TO15(-762305), .W51TO16(466919), .W51TO17(630397), .W51TO18(62550), .W51TO19(-782030), .W51TO20(480471), .W51TO21(531114), .W51TO22(714930), .W51TO23(214978), .W51TO24(564330), .W51TO25(-180511), .W51TO26(889108), .W51TO27(-525025), .W51TO28(-408829), .W51TO29(-629738), .W51TO30(786171), .W51TO31(-484699), .W51TO32(132062), .W51TO33(479120), .W51TO34(870277), .W51TO35(309039), .W51TO36(318411), .W51TO37(-943537), .W51TO38(358737), .W51TO39(270953), .W51TO40(-695779), .W51TO41(531332), .W51TO42(-438819), .W51TO43(-47024), .W51TO44(-464434), .W51TO45(771376), .W51TO46(918354), .W51TO47(-511258), .W51TO48(921291), .W51TO49(-39680), .W51TO50(351891), .W51TO51(714657), .W51TO52(-731703), .W51TO53(-217751), .W51TO54(-256435), .W51TO55(899454), .W51TO56(-475020), .W51TO57(813505), .W51TO58(-905367), .W51TO59(-929366), .W51TO60(534799), .W51TO61(-210946), .W51TO62(-58108), .W51TO63(247552), .W52TO0(727483), .W52TO1(919508), .W52TO2(-755293), .W52TO3(-767797), .W52TO4(-887904), .W52TO5(-586797), .W52TO6(955630), .W52TO7(-607472), .W52TO8(243539), .W52TO9(-497568), .W52TO10(-53068), .W52TO11(-396134), .W52TO12(293811), .W52TO13(845134), .W52TO14(-233068), .W52TO15(570099), .W52TO16(237563), .W52TO17(-323672), .W52TO18(762953), .W52TO19(-846433), .W52TO20(45174), .W52TO21(-545823), .W52TO22(-446857), .W52TO23(343450), .W52TO24(700008), .W52TO25(748698), .W52TO26(787291), .W52TO27(952453), .W52TO28(458350), .W52TO29(-598832), .W52TO30(-749345), .W52TO31(55661), .W52TO32(233756), .W52TO33(65768), .W52TO34(911193), .W52TO35(746299), .W52TO36(-559436), .W52TO37(35692), .W52TO38(389314), .W52TO39(472231), .W52TO40(84956), .W52TO41(-279116), .W52TO42(819862), .W52TO43(419784), .W52TO44(988114), .W52TO45(-278879), .W52TO46(504224), .W52TO47(-770202), .W52TO48(-968892), .W52TO49(-611932), .W52TO50(-683595), .W52TO51(-276211), .W52TO52(345552), .W52TO53(81887), .W52TO54(-594515), .W52TO55(-33674), .W52TO56(521251), .W52TO57(782847), .W52TO58(745839), .W52TO59(-527886), .W52TO60(-161279), .W52TO61(485312), .W52TO62(777873), .W52TO63(175905), .W53TO0(307103), .W53TO1(387120), .W53TO2(-664929), .W53TO3(-334403), .W53TO4(-408014), .W53TO5(-989619), .W53TO6(986839), .W53TO7(218763), .W53TO8(916880), .W53TO9(923897), .W53TO10(-745751), .W53TO11(263133), .W53TO12(162427), .W53TO13(-72666), .W53TO14(131164), .W53TO15(72028), .W53TO16(-393051), .W53TO17(906427), .W53TO18(-949545), .W53TO19(822303), .W53TO20(110852), .W53TO21(609601), .W53TO22(-831445), .W53TO23(-863332), .W53TO24(-976660), .W53TO25(265499), .W53TO26(564027), .W53TO27(799181), .W53TO28(-156030), .W53TO29(338993), .W53TO30(15604), .W53TO31(235465), .W53TO32(-147992), .W53TO33(-458211), .W53TO34(899976), .W53TO35(-179105), .W53TO36(-345211), .W53TO37(-195260), .W53TO38(520949), .W53TO39(976986), .W53TO40(651693), .W53TO41(913892), .W53TO42(1770), .W53TO43(-981914), .W53TO44(-41883), .W53TO45(-946589), .W53TO46(879442), .W53TO47(-49194), .W53TO48(904250), .W53TO49(312900), .W53TO50(962040), .W53TO51(-717470), .W53TO52(566855), .W53TO53(713951), .W53TO54(-605412), .W53TO55(523555), .W53TO56(-758380), .W53TO57(98353), .W53TO58(-188818), .W53TO59(-402580), .W53TO60(703539), .W53TO61(758717), .W53TO62(318019), .W53TO63(-179380), .W54TO0(-719455), .W54TO1(-408303), .W54TO2(853917), .W54TO3(-94172), .W54TO4(-53138), .W54TO5(619099), .W54TO6(-563717), .W54TO7(289566), .W54TO8(875957), .W54TO9(-43664), .W54TO10(572430), .W54TO11(-315167), .W54TO12(-6578), .W54TO13(780541), .W54TO14(-566304), .W54TO15(981364), .W54TO16(-822129), .W54TO17(577449), .W54TO18(680682), .W54TO19(355312), .W54TO20(925109), .W54TO21(-41318), .W54TO22(435835), .W54TO23(362226), .W54TO24(-689299), .W54TO25(804895), .W54TO26(516186), .W54TO27(858877), .W54TO28(243262), .W54TO29(-946960), .W54TO30(265227), .W54TO31(-319447), .W54TO32(190680), .W54TO33(282724), .W54TO34(-309245), .W54TO35(417756), .W54TO36(-669804), .W54TO37(400400), .W54TO38(221972), .W54TO39(-664201), .W54TO40(757702), .W54TO41(-266097), .W54TO42(922104), .W54TO43(-333798), .W54TO44(-432275), .W54TO45(-399837), .W54TO46(806077), .W54TO47(-558808), .W54TO48(-976208), .W54TO49(334046), .W54TO50(538577), .W54TO51(190351), .W54TO52(625940), .W54TO53(149915), .W54TO54(-238437), .W54TO55(-767092), .W54TO56(16006), .W54TO57(536858), .W54TO58(-950436), .W54TO59(569516), .W54TO60(264598), .W54TO61(-592973), .W54TO62(-632787), .W54TO63(431591), .W55TO0(623946), .W55TO1(-857882), .W55TO2(986156), .W55TO3(505530), .W55TO4(129425), .W55TO5(-409754), .W55TO6(-289022), .W55TO7(-176510), .W55TO8(-270182), .W55TO9(-15555), .W55TO10(352996), .W55TO11(839369), .W55TO12(586342), .W55TO13(-71607), .W55TO14(413019), .W55TO15(879194), .W55TO16(841671), .W55TO17(189176), .W55TO18(905157), .W55TO19(395028), .W55TO20(590980), .W55TO21(148966), .W55TO22(132198), .W55TO23(584232), .W55TO24(971845), .W55TO25(-916680), .W55TO26(-107710), .W55TO27(-928142), .W55TO28(821365), .W55TO29(132986), .W55TO30(-844977), .W55TO31(-391318), .W55TO32(-390076), .W55TO33(966052), .W55TO34(-254194), .W55TO35(209338), .W55TO36(-803750), .W55TO37(-124245), .W55TO38(-285981), .W55TO39(-325453), .W55TO40(-858086), .W55TO41(973025), .W55TO42(-428251), .W55TO43(520706), .W55TO44(-30185), .W55TO45(-968837), .W55TO46(-765201), .W55TO47(-542712), .W55TO48(-461894), .W55TO49(699275), .W55TO50(-502508), .W55TO51(300295), .W55TO52(591879), .W55TO53(-470369), .W55TO54(-270416), .W55TO55(90114), .W55TO56(801622), .W55TO57(373885), .W55TO58(-889490), .W55TO59(975273), .W55TO60(-931322), .W55TO61(655175), .W55TO62(-771769), .W55TO63(723320), .W56TO0(-458186), .W56TO1(-419200), .W56TO2(-590937), .W56TO3(904648), .W56TO4(-966842), .W56TO5(556679), .W56TO6(273808), .W56TO7(740361), .W56TO8(35685), .W56TO9(-40668), .W56TO10(-972735), .W56TO11(294708), .W56TO12(160961), .W56TO13(222996), .W56TO14(-397084), .W56TO15(716595), .W56TO16(13297), .W56TO17(135666), .W56TO18(711447), .W56TO19(-365153), .W56TO20(115143), .W56TO21(-463681), .W56TO22(-287249), .W56TO23(595575), .W56TO24(363730), .W56TO25(-914508), .W56TO26(-14631), .W56TO27(-877455), .W56TO28(-591747), .W56TO29(200656), .W56TO30(-114568), .W56TO31(-487099), .W56TO32(41156), .W56TO33(-235206), .W56TO34(-498029), .W56TO35(191645), .W56TO36(770742), .W56TO37(-505621), .W56TO38(-425321), .W56TO39(-602852), .W56TO40(-599526), .W56TO41(-195997), .W56TO42(893422), .W56TO43(-605582), .W56TO44(-884561), .W56TO45(-83344), .W56TO46(793019), .W56TO47(-812664), .W56TO48(172905), .W56TO49(962328), .W56TO50(-608341), .W56TO51(407475), .W56TO52(-438809), .W56TO53(746381), .W56TO54(352258), .W56TO55(397677), .W56TO56(301868), .W56TO57(-986114), .W56TO58(791160), .W56TO59(925425), .W56TO60(549616), .W56TO61(343606), .W56TO62(45108), .W56TO63(482881), .W57TO0(-805058), .W57TO1(-967544), .W57TO2(960549), .W57TO3(-67586), .W57TO4(-607109), .W57TO5(522401), .W57TO6(-982083), .W57TO7(-876739), .W57TO8(98884), .W57TO9(874101), .W57TO10(739149), .W57TO11(811630), .W57TO12(-625026), .W57TO13(920307), .W57TO14(-813767), .W57TO15(-736312), .W57TO16(354321), .W57TO17(903538), .W57TO18(49368), .W57TO19(-104341), .W57TO20(-486032), .W57TO21(962726), .W57TO22(129082), .W57TO23(-839962), .W57TO24(-129195), .W57TO25(57651), .W57TO26(-994808), .W57TO27(-85249), .W57TO28(410518), .W57TO29(32060), .W57TO30(-430889), .W57TO31(399206), .W57TO32(808393), .W57TO33(947289), .W57TO34(-874093), .W57TO35(98089), .W57TO36(88705), .W57TO37(681192), .W57TO38(661693), .W57TO39(-10381), .W57TO40(-438673), .W57TO41(585344), .W57TO42(345222), .W57TO43(-251018), .W57TO44(-890357), .W57TO45(892279), .W57TO46(-299713), .W57TO47(62249), .W57TO48(-146684), .W57TO49(60170), .W57TO50(-837052), .W57TO51(-319601), .W57TO52(-948200), .W57TO53(-662060), .W57TO54(286681), .W57TO55(883490), .W57TO56(343633), .W57TO57(-38976), .W57TO58(789716), .W57TO59(-27415), .W57TO60(-743470), .W57TO61(-574993), .W57TO62(177728), .W57TO63(-113269), .W58TO0(-621980), .W58TO1(392010), .W58TO2(-286820), .W58TO3(-13051), .W58TO4(656768), .W58TO5(271665), .W58TO6(728809), .W58TO7(-314563), .W58TO8(840132), .W58TO9(-623171), .W58TO10(-394102), .W58TO11(-691039), .W58TO12(-585251), .W58TO13(-305998), .W58TO14(-530380), .W58TO15(-163167), .W58TO16(619814), .W58TO17(-928150), .W58TO18(-201591), .W58TO19(-989805), .W58TO20(793125), .W58TO21(272485), .W58TO22(149188), .W58TO23(639453), .W58TO24(945439), .W58TO25(849025), .W58TO26(-42536), .W58TO27(635175), .W58TO28(-59833), .W58TO29(-65671), .W58TO30(437016), .W58TO31(509985), .W58TO32(719947), .W58TO33(-62848), .W58TO34(296963), .W58TO35(131819), .W58TO36(474883), .W58TO37(69186), .W58TO38(198485), .W58TO39(-728173), .W58TO40(-68283), .W58TO41(-208974), .W58TO42(-723225), .W58TO43(-207198), .W58TO44(226512), .W58TO45(-732874), .W58TO46(741048), .W58TO47(90224), .W58TO48(311409), .W58TO49(-88458), .W58TO50(307965), .W58TO51(-748073), .W58TO52(-546485), .W58TO53(-757516), .W58TO54(373474), .W58TO55(-503166), .W58TO56(-89217), .W58TO57(-179222), .W58TO58(994161), .W58TO59(749979), .W58TO60(-419980), .W58TO61(804937), .W58TO62(287307), .W58TO63(260561), .W59TO0(-322822), .W59TO1(782831), .W59TO2(504572), .W59TO3(-760797), .W59TO4(267880), .W59TO5(-835336), .W59TO6(651997), .W59TO7(889214), .W59TO8(-792491), .W59TO9(-711103), .W59TO10(-433696), .W59TO11(-224279), .W59TO12(-545378), .W59TO13(645305), .W59TO14(-172844), .W59TO15(932138), .W59TO16(-860935), .W59TO17(974024), .W59TO18(259465), .W59TO19(-297972), .W59TO20(-660617), .W59TO21(-89230), .W59TO22(-83903), .W59TO23(409075), .W59TO24(836347), .W59TO25(-747566), .W59TO26(-93359), .W59TO27(328956), .W59TO28(140187), .W59TO29(201760), .W59TO30(-776451), .W59TO31(969829), .W59TO32(-25419), .W59TO33(-785945), .W59TO34(-769258), .W59TO35(205618), .W59TO36(-888571), .W59TO37(219562), .W59TO38(-811883), .W59TO39(754222), .W59TO40(458900), .W59TO41(558320), .W59TO42(-297393), .W59TO43(403620), .W59TO44(112659), .W59TO45(-73876), .W59TO46(370397), .W59TO47(-879055), .W59TO48(-116417), .W59TO49(-516643), .W59TO50(-825044), .W59TO51(-496265), .W59TO52(-999115), .W59TO53(986240), .W59TO54(103552), .W59TO55(510658), .W59TO56(-872534), .W59TO57(-707698), .W59TO58(467093), .W59TO59(648973), .W59TO60(640846), .W59TO61(-81051), .W59TO62(-769467), .W59TO63(398764), .W60TO0(-84523), .W60TO1(-217668), .W60TO2(-732840), .W60TO3(-818774), .W60TO4(449085), .W60TO5(576416), .W60TO6(606408), .W60TO7(888086), .W60TO8(-476667), .W60TO9(-817534), .W60TO10(518668), .W60TO11(-305080), .W60TO12(-985064), .W60TO13(-419473), .W60TO14(280338), .W60TO15(-568140), .W60TO16(-195659), .W60TO17(-977760), .W60TO18(-952750), .W60TO19(490576), .W60TO20(191587), .W60TO21(344331), .W60TO22(-469255), .W60TO23(-528873), .W60TO24(527539), .W60TO25(-344893), .W60TO26(763487), .W60TO27(-729357), .W60TO28(-971312), .W60TO29(-34850), .W60TO30(779663), .W60TO31(386129), .W60TO32(-670457), .W60TO33(-751356), .W60TO34(511284), .W60TO35(124897), .W60TO36(72049), .W60TO37(-927148), .W60TO38(167928), .W60TO39(-451190), .W60TO40(710081), .W60TO41(-638563), .W60TO42(-777515), .W60TO43(-665844), .W60TO44(722084), .W60TO45(435754), .W60TO46(150361), .W60TO47(-222390), .W60TO48(-767134), .W60TO49(139596), .W60TO50(-261342), .W60TO51(-792581), .W60TO52(-495129), .W60TO53(-800148), .W60TO54(-830996), .W60TO55(-310906), .W60TO56(954998), .W60TO57(111550), .W60TO58(484706), .W60TO59(651803), .W60TO60(-204622), .W60TO61(650608), .W60TO62(11439), .W60TO63(823526), .W61TO0(529136), .W61TO1(651844), .W61TO2(360508), .W61TO3(669257), .W61TO4(719915), .W61TO5(169789), .W61TO6(619238), .W61TO7(741205), .W61TO8(546072), .W61TO9(821185), .W61TO10(-586478), .W61TO11(219177), .W61TO12(-994756), .W61TO13(73454), .W61TO14(635046), .W61TO15(592907), .W61TO16(-160569), .W61TO17(-235346), .W61TO18(706732), .W61TO19(-157971), .W61TO20(331281), .W61TO21(602249), .W61TO22(-540163), .W61TO23(248330), .W61TO24(-565606), .W61TO25(-92926), .W61TO26(47955), .W61TO27(904392), .W61TO28(938351), .W61TO29(-494127), .W61TO30(409092), .W61TO31(621956), .W61TO32(-624351), .W61TO33(513074), .W61TO34(-77713), .W61TO35(-20437), .W61TO36(306338), .W61TO37(465928), .W61TO38(-505561), .W61TO39(-498169), .W61TO40(925537), .W61TO41(864654), .W61TO42(437946), .W61TO43(-106871), .W61TO44(-203647), .W61TO45(68322), .W61TO46(-990724), .W61TO47(372292), .W61TO48(321563), .W61TO49(814391), .W61TO50(-727258), .W61TO51(-657303), .W61TO52(-710014), .W61TO53(650772), .W61TO54(39030), .W61TO55(979146), .W61TO56(-578826), .W61TO57(236872), .W61TO58(464900), .W61TO59(-234101), .W61TO60(-877075), .W61TO61(-193068), .W61TO62(-558799), .W61TO63(-34520), .W62TO0(-327485), .W62TO1(492988), .W62TO2(642860), .W62TO3(706358), .W62TO4(485921), .W62TO5(122670), .W62TO6(664372), .W62TO7(431215), .W62TO8(234064), .W62TO9(938213), .W62TO10(-918758), .W62TO11(-451403), .W62TO12(589133), .W62TO13(-766234), .W62TO14(-641377), .W62TO15(672126), .W62TO16(-320640), .W62TO17(-385332), .W62TO18(-102538), .W62TO19(-211570), .W62TO20(931718), .W62TO21(-660876), .W62TO22(-701041), .W62TO23(-963210), .W62TO24(624075), .W62TO25(-711640), .W62TO26(-947746), .W62TO27(321956), .W62TO28(-760731), .W62TO29(-723638), .W62TO30(-103513), .W62TO31(-155469), .W62TO32(242428), .W62TO33(-453478), .W62TO34(935296), .W62TO35(-540001), .W62TO36(-212387), .W62TO37(-817128), .W62TO38(-665000), .W62TO39(-936612), .W62TO40(313212), .W62TO41(-92063), .W62TO42(599595), .W62TO43(-217719), .W62TO44(-985911), .W62TO45(606547), .W62TO46(-947055), .W62TO47(-366412), .W62TO48(597368), .W62TO49(196822), .W62TO50(720071), .W62TO51(478102), .W62TO52(-898315), .W62TO53(272531), .W62TO54(-369712), .W62TO55(822274), .W62TO56(-88681), .W62TO57(768471), .W62TO58(-493920), .W62TO59(54588), .W62TO60(-912770), .W62TO61(-595498), .W62TO62(947248), .W62TO63(-948537), .W63TO0(846112), .W63TO1(699823), .W63TO2(-502420), .W63TO3(-998592), .W63TO4(473896), .W63TO5(731501), .W63TO6(-619070), .W63TO7(951296), .W63TO8(876729), .W63TO9(541429), .W63TO10(-447574), .W63TO11(725942), .W63TO12(324861), .W63TO13(768422), .W63TO14(18706), .W63TO15(708900), .W63TO16(286402), .W63TO17(-784284), .W63TO18(-536046), .W63TO19(6707), .W63TO20(-401131), .W63TO21(129267), .W63TO22(-724128), .W63TO23(-289945), .W63TO24(501504), .W63TO25(474720), .W63TO26(250705), .W63TO27(-469645), .W63TO28(-881137), .W63TO29(-124528), .W63TO30(732360), .W63TO31(646458), .W63TO32(721745), .W63TO33(-407522), .W63TO34(869331), .W63TO35(-190111), .W63TO36(-977438), .W63TO37(-326028), .W63TO38(422747), .W63TO39(-722184), .W63TO40(803311), .W63TO41(533705), .W63TO42(664263), .W63TO43(540630), .W63TO44(-42154), .W63TO45(633693), .W63TO46(-951284), .W63TO47(-160793), .W63TO48(284140), .W63TO49(963287), .W63TO50(-972793), .W63TO51(-335716), .W63TO52(121153), .W63TO53(93008), .W63TO54(-96388), .W63TO55(-253089), .W63TO56(960999), .W63TO57(796107), .W63TO58(-493484), .W63TO59(-836392), .W63TO60(609971), .W63TO61(624649), .W63TO62(-592088), .W63TO63(313160), .W64TO0(-251528), .W64TO1(-842571), .W64TO2(796481), .W64TO3(-963446), .W64TO4(302467), .W64TO5(491966), .W64TO6(-623231), .W64TO7(796468), .W64TO8(557592), .W64TO9(548681), .W64TO10(-530714), .W64TO11(-729727), .W64TO12(991602), .W64TO13(612354), .W64TO14(-255413), .W64TO15(-751645), .W64TO16(708247), .W64TO17(-835445), .W64TO18(-666725), .W64TO19(-754882), .W64TO20(-601319), .W64TO21(-73275), .W64TO22(-664087), .W64TO23(810828), .W64TO24(-173320), .W64TO25(-199222), .W64TO26(-509822), .W64TO27(33220), .W64TO28(29290), .W64TO29(931938), .W64TO30(677731), .W64TO31(544310), .W64TO32(-346977), .W64TO33(569614), .W64TO34(161950), .W64TO35(-58199), .W64TO36(-429742), .W64TO37(621776), .W64TO38(433984), .W64TO39(237583), .W64TO40(-916969), .W64TO41(290548), .W64TO42(302206), .W64TO43(-724057), .W64TO44(-503723), .W64TO45(783758), .W64TO46(989933), .W64TO47(56120), .W64TO48(-780769), .W64TO49(-102667), .W64TO50(727677), .W64TO51(214598), .W64TO52(23844), .W64TO53(889952), .W64TO54(-526709), .W64TO55(-938643), .W64TO56(-830338), .W64TO57(-932592), .W64TO58(-986098), .W64TO59(-672417), .W64TO60(171935), .W64TO61(231598), .W64TO62(-187399), .W64TO63(-692766)) layer0(.clk(clk), .rst(rst), .in0(in0), .in1(in1), .in2(in2), .in3(in3), .in4(in4), .in5(in5), .in6(in6), .in7(in7), .in8(in8), .in9(in9), .in10(in10), .in11(in11), .in12(in12), .in13(in13), .in14(in14), .in15(in15), .in16(in16), .in17(in17), .in18(in18), .in19(in19), .in20(in20), .in21(in21), .in22(in22), .in23(in23), .in24(in24), .in25(in25), .in26(in26), .in27(in27), .in28(in28), .in29(in29), .in30(in30), .in31(in31), .in32(in32), .in33(in33), .in34(in34), .in35(in35), .in36(in36), .in37(in37), .in38(in38), .in39(in39), .in40(in40), .in41(in41), .in42(in42), .in43(in43), .in44(in44), .in45(in45), .in46(in46), .in47(in47), .in48(in48), .in49(in49), .in50(in50), .in51(in51), .in52(in52), .in53(in53), .in54(in54), .in55(in55), .in56(in56), .in57(in57), .in58(in58), .in59(in59), .in60(in60), .in61(in61), .in62(in62), .in63(in63), .in64(in64), .out0(con0[0]), .out1(con0[1]), .out2(con0[2]), .out3(con0[3]), .out4(con0[4]), .out5(con0[5]), .out6(con0[6]), .out7(con0[7]), .out8(con0[8]), .out9(con0[9]), .out10(con0[10]), .out11(con0[11]), .out12(con0[12]), .out13(con0[13]), .out14(con0[14]), .out15(con0[15]), .out16(con0[16]), .out17(con0[17]), .out18(con0[18]), .out19(con0[19]), .out20(con0[20]), .out21(con0[21]), .out22(con0[22]), .out23(con0[23]), .out24(con0[24]), .out25(con0[25]), .out26(con0[26]), .out27(con0[27]), .out28(con0[28]), .out29(con0[29]), .out30(con0[30]), .out31(con0[31]), .out32(con0[32]), .out33(con0[33]), .out34(con0[34]), .out35(con0[35]), .out36(con0[36]), .out37(con0[37]), .out38(con0[38]), .out39(con0[39]), .out40(con0[40]), .out41(con0[41]), .out42(con0[42]), .out43(con0[43]), .out44(con0[44]), .out45(con0[45]), .out46(con0[46]), .out47(con0[47]), .out48(con0[48]), .out49(con0[49]), .out50(con0[50]), .out51(con0[51]), .out52(con0[52]), .out53(con0[53]), .out54(con0[54]), .out55(con0[55]), .out56(con0[56]), .out57(con0[57]), .out58(con0[58]), .out59(con0[59]), .out60(con0[60]), .out61(con0[61]), .out62(con0[62]), .out63(con0[63]));
layer64in1out #(.BIAS0(-917974), .W0TO0(970580), .W1TO0(-583174), .W2TO0(-108499), .W3TO0(-947074), .W4TO0(10114), .W5TO0(-181164), .W6TO0(-751155), .W7TO0(-765588), .W8TO0(916346), .W9TO0(973126), .W10TO0(779388), .W11TO0(-737647), .W12TO0(190585), .W13TO0(-446431), .W14TO0(310802), .W15TO0(-970128), .W16TO0(-173047), .W17TO0(-606779), .W18TO0(-20357), .W19TO0(73388), .W20TO0(669226), .W21TO0(-147587), .W22TO0(865480), .W23TO0(-846169), .W24TO0(-158879), .W25TO0(836912), .W26TO0(-714310), .W27TO0(-403376), .W28TO0(-159168), .W29TO0(39759), .W30TO0(-371807), .W31TO0(576669), .W32TO0(-86168), .W33TO0(-501811), .W34TO0(-221142), .W35TO0(545212), .W36TO0(-483003), .W37TO0(-271982), .W38TO0(-342895), .W39TO0(-641355), .W40TO0(766762), .W41TO0(-507131), .W42TO0(-804702), .W43TO0(215568), .W44TO0(992350), .W45TO0(274023), .W46TO0(550710), .W47TO0(563961), .W48TO0(-579716), .W49TO0(-632364), .W50TO0(141114), .W51TO0(-562972), .W52TO0(850542), .W53TO0(207935), .W54TO0(111886), .W55TO0(-139913), .W56TO0(-533575), .W57TO0(304183), .W58TO0(957052), .W59TO0(219720), .W60TO0(952251), .W61TO0(-95299), .W62TO0(-155802), .W63TO0(20059)) layer1(.clk(clk), .rst(rst), .in0(con0[0]), .in1(con0[1]), .in2(con0[2]), .in3(con0[3]), .in4(con0[4]), .in5(con0[5]), .in6(con0[6]), .in7(con0[7]), .in8(con0[8]), .in9(con0[9]), .in10(con0[10]), .in11(con0[11]), .in12(con0[12]), .in13(con0[13]), .in14(con0[14]), .in15(con0[15]), .in16(con0[16]), .in17(con0[17]), .in18(con0[18]), .in19(con0[19]), .in20(con0[20]), .in21(con0[21]), .in22(con0[22]), .in23(con0[23]), .in24(con0[24]), .in25(con0[25]), .in26(con0[26]), .in27(con0[27]), .in28(con0[28]), .in29(con0[29]), .in30(con0[30]), .in31(con0[31]), .in32(con0[32]), .in33(con0[33]), .in34(con0[34]), .in35(con0[35]), .in36(con0[36]), .in37(con0[37]), .in38(con0[38]), .in39(con0[39]), .in40(con0[40]), .in41(con0[41]), .in42(con0[42]), .in43(con0[43]), .in44(con0[44]), .in45(con0[45]), .in46(con0[46]), .in47(con0[47]), .in48(con0[48]), .in49(con0[49]), .in50(con0[50]), .in51(con0[51]), .in52(con0[52]), .in53(con0[53]), .in54(con0[54]), .in55(con0[55]), .in56(con0[56]), .in57(con0[57]), .in58(con0[58]), .in59(con0[59]), .in60(con0[60]), .in61(con0[61]), .in62(con0[62]), .in63(con0[63]), .out0(out0));

endmodule

`define assert_close(expected, got, eps) \
if ((expected > got && expected > got + eps) || (expected < got && expected + eps < got)) begin \
    $display("TEST FAILED in %m: got %d, expected %d", got, expected); \
end

module example_tb;
logic clk;
logic rst;

reg signed [63:0] net_in0, net_in1, net_in2, net_in3, net_in4, net_in5, net_in6, net_in7, net_in8, net_in9, net_in10, net_in11, net_in12, net_in13, net_in14, net_in15, net_in16, net_in17, net_in18, net_in19, net_in20, net_in21, net_in22, net_in23, net_in24, net_in25, net_in26, net_in27, net_in28, net_in29, net_in30, net_in31, net_in32, net_in33, net_in34, net_in35, net_in36, net_in37, net_in38, net_in39, net_in40, net_in41, net_in42, net_in43, net_in44, net_in45, net_in46, net_in47, net_in48, net_in49, net_in50, net_in51, net_in52, net_in53, net_in54, net_in55, net_in56, net_in57, net_in58, net_in59, net_in60, net_in61, net_in62, net_in63, net_in64;

wire signed [63:0] net_out0;

network net(.clk(clk), .rst(rst), .in0(net_in0), .in1(net_in1), .in2(net_in2), .in3(net_in3), .in4(net_in4), .in5(net_in5), .in6(net_in6), .in7(net_in7), .in8(net_in8), .in9(net_in9), .in10(net_in10), .in11(net_in11), .in12(net_in12), .in13(net_in13), .in14(net_in14), .in15(net_in15), .in16(net_in16), .in17(net_in17), .in18(net_in18), .in19(net_in19), .in20(net_in20), .in21(net_in21), .in22(net_in22), .in23(net_in23), .in24(net_in24), .in25(net_in25), .in26(net_in26), .in27(net_in27), .in28(net_in28), .in29(net_in29), .in30(net_in30), .in31(net_in31), .in32(net_in32), .in33(net_in33), .in34(net_in34), .in35(net_in35), .in36(net_in36), .in37(net_in37), .in38(net_in38), .in39(net_in39), .in40(net_in40), .in41(net_in41), .in42(net_in42), .in43(net_in43), .in44(net_in44), .in45(net_in45), .in46(net_in46), .in47(net_in47), .in48(net_in48), .in49(net_in49), .in50(net_in50), .in51(net_in51), .in52(net_in52), .in53(net_in53), .in54(net_in54), .in55(net_in55), .in56(net_in56), .in57(net_in57), .in58(net_in58), .in59(net_in59), .in60(net_in60), .in61(net_in61), .in62(net_in62), .in63(net_in63), .in64(net_in64), .out0(net_out0));

task test;
input signed [63:0] in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31, in32, in33, in34, in35, in36, in37, in38, in39, in40, in41, in42, in43, in44, in45, in46, in47, in48, in49, in50, in51, in52, in53, in54, in55, in56, in57, in58, in59, in60, in61, in62, in63, in64, out0;
begin
    net_in0 = in0;
    net_in1 = in1;
    net_in2 = in2;
    net_in3 = in3;
    net_in4 = in4;
    net_in5 = in5;
    net_in6 = in6;
    net_in7 = in7;
    net_in8 = in8;
    net_in9 = in9;
    net_in10 = in10;
    net_in11 = in11;
    net_in12 = in12;
    net_in13 = in13;
    net_in14 = in14;
    net_in15 = in15;
    net_in16 = in16;
    net_in17 = in17;
    net_in18 = in18;
    net_in19 = in19;
    net_in20 = in20;
    net_in21 = in21;
    net_in22 = in22;
    net_in23 = in23;
    net_in24 = in24;
    net_in25 = in25;
    net_in26 = in26;
    net_in27 = in27;
    net_in28 = in28;
    net_in29 = in29;
    net_in30 = in30;
    net_in31 = in31;
    net_in32 = in32;
    net_in33 = in33;
    net_in34 = in34;
    net_in35 = in35;
    net_in36 = in36;
    net_in37 = in37;
    net_in38 = in38;
    net_in39 = in39;
    net_in40 = in40;
    net_in41 = in41;
    net_in42 = in42;
    net_in43 = in43;
    net_in44 = in44;
    net_in45 = in45;
    net_in46 = in46;
    net_in47 = in47;
    net_in48 = in48;
    net_in49 = in49;
    net_in50 = in50;
    net_in51 = in51;
    net_in52 = in52;
    net_in53 = in53;
    net_in54 = in54;
    net_in55 = in55;
    net_in56 = in56;
    net_in57 = in57;
    net_in58 = in58;
    net_in59 = in59;
    net_in60 = in60;
    net_in61 = in61;
    net_in62 = in62;
    net_in63 = in63;
    net_in64 = in64;
    #10000000ns
    `assert_close(out0, net_out0, 10000);
end
endtask

initial
begin
    $dumpfile("waves.vcd");
    $dumpvars;
    test(0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 215436);
    $display("Test0 completed");
    test(1000000, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 160313);
    $display("Test1 completed");
    test(0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 626831);
    $display("Test2 completed");
    test(0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 58821);
    $display("Test3 completed");
    test(1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 0, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 57350);
    $display("Test4 completed");
    test(0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 0, 74383);
    $display("Test5 completed");
    test(0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 597126);
    $display("Test6 completed");
    test(1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 120165);
    $display("Test7 completed");
    test(1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 130793);
    $display("Test8 completed");
    test(0, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 66971);
    $display("Test9 completed");
    test(1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 72279);
    $display("Test10 completed");
    test(0, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 0, 58484);
    $display("Test11 completed");
    test(1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 292957);
    $display("Test12 completed");
    test(1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 81472);
    $display("Test13 completed");
    test(0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 288623);
    $display("Test14 completed");
    test(0, 0, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 75673);
    $display("Test15 completed");
    test(0, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 126353);
    $display("Test16 completed");
    test(0, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 80675);
    $display("Test17 completed");
    test(0, 0, 0, 1000000, 0, 1000000, 0, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 290242);
    $display("Test18 completed");
    test(1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 115135);
    $display("Test19 completed");
    test(1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 1000000, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 0, 136485);
    $display("Test20 completed");
    test(0, 0, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 151643);
    $display("Test21 completed");
    test(0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 324266);
    $display("Test22 completed");
    test(1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 0, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 522330);
    $display("Test23 completed");
    test(1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 663980);
    $display("Test24 completed");
    test(0, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 501861);
    $display("Test25 completed");
    test(1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 0, 179144);
    $display("Test26 completed");
    test(1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 0, 302377);
    $display("Test27 completed");
    test(0, 1000000, 0, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 142492);
    $display("Test28 completed");
    test(0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 465726);
    $display("Test29 completed");
    test(0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 0, 77812);
    $display("Test30 completed");
    test(1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 0, 0, 482046);
    $display("Test31 completed");
    test(0, 1000000, 0, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 163454);
    $display("Test32 completed");
    test(0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 217831);
    $display("Test33 completed");
    test(0, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 0, 0, 1000000, 228690);
    $display("Test34 completed");
    test(0, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 0, 1000000, 0, 1000000, 331620);
    $display("Test35 completed");
    test(0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 0, 0, 98556);
    $display("Test36 completed");
    test(1000000, 0, 0, 1000000, 0, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 164029);
    $display("Test37 completed");
    test(1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 107753);
    $display("Test38 completed");
    test(1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 254192);
    $display("Test39 completed");
    test(1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 0, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 358735);
    $display("Test40 completed");
    test(0, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 69907);
    $display("Test41 completed");
    test(1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 130326);
    $display("Test42 completed");
    test(0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 0, 195178);
    $display("Test43 completed");
    test(0, 1000000, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 347904);
    $display("Test44 completed");
    test(1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 156171);
    $display("Test45 completed");
    test(1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 9428);
    $display("Test46 completed");
    test(0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 0, 85202);
    $display("Test47 completed");
    test(0, 1000000, 1000000, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 138497);
    $display("Test48 completed");
    test(0, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 51400);
    $display("Test49 completed");
    test(0, 0, 0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 77796);
    $display("Test50 completed");
    test(1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 157204);
    $display("Test51 completed");
    test(0, 0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 0, 185880);
    $display("Test52 completed");
    test(1000000, 0, 0, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 63961);
    $display("Test53 completed");
    test(1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 188324);
    $display("Test54 completed");
    test(1000000, 1000000, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 210420);
    $display("Test55 completed");
    test(0, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 46748);
    $display("Test56 completed");
    test(0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 53982);
    $display("Test57 completed");
    test(0, 1000000, 1000000, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 433027);
    $display("Test58 completed");
    test(0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 778035);
    $display("Test59 completed");
    test(1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 331354);
    $display("Test60 completed");
    test(0, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 151779);
    $display("Test61 completed");
    test(1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 0, 1000000, 1000000, 0, 0, 0, 386637);
    $display("Test62 completed");
    test(1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 0, 0, 181707);
    $display("Test63 completed");
    test(1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 238732);
    $display("Test64 completed");
    test(0, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 267568);
    $display("Test65 completed");
    test(1000000, 0, 0, 1000000, 0, 0, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 683365);
    $display("Test66 completed");
    test(1000000, 0, 0, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 1000000, 1000000, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 1000000, 58531);
    $display("Test67 completed");
    test(0, 0, 0, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 114024);
    $display("Test68 completed");
    test(1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 39204);
    $display("Test69 completed");
    test(0, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 99181);
    $display("Test70 completed");
    test(0, 1000000, 0, 0, 0, 0, 0, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 785361);
    $display("Test71 completed");
    test(0, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 114575);
    $display("Test72 completed");
    test(0, 0, 1000000, 0, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 143477);
    $display("Test73 completed");
    test(0, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 705264);
    $display("Test74 completed");
    test(1000000, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 178926);
    $display("Test75 completed");
    test(1000000, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 196422);
    $display("Test76 completed");
    test(0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 227623);
    $display("Test77 completed");
    test(1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 0, 60484);
    $display("Test78 completed");
    test(1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 73221);
    $display("Test79 completed");
    test(1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 510136);
    $display("Test80 completed");
    test(0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 256667);
    $display("Test81 completed");
    test(1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 40584);
    $display("Test82 completed");
    test(0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 248281);
    $display("Test83 completed");
    test(0, 1000000, 0, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 0, 1000000, 0, 0, 353515);
    $display("Test84 completed");
    test(0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 165883);
    $display("Test85 completed");
    test(0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 80196);
    $display("Test86 completed");
    test(1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 271233);
    $display("Test87 completed");
    test(0, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 210973);
    $display("Test88 completed");
    test(0, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 675583);
    $display("Test89 completed");
    test(1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 166083);
    $display("Test90 completed");
    test(0, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 61353);
    $display("Test91 completed");
    test(0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 391060);
    $display("Test92 completed");
    test(0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 60420);
    $display("Test93 completed");
    test(1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 0, 1000000, 0, 0, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 71807);
    $display("Test94 completed");
    test(1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 0, 101939);
    $display("Test95 completed");
    test(0, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 49610);
    $display("Test96 completed");
    test(1000000, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 0, 1000000, 0, 0, 1000000, 74273);
    $display("Test97 completed");
    test(1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 1000000, 0, 1000000, 0, 1000000, 1000000, 0, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 1000000, 0, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 31017);
    $display("Test98 completed");
    test(0, 1000000, 0, 1000000, 0, 0, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 1000000, 0, 1000000, 1000000, 0, 0, 1000000, 1000000, 0, 0, 1000000, 0, 0, 1000000, 1000000, 0, 0, 0, 0, 0, 1000000, 1000000, 1000000, 1000000, 0, 0, 0, 0, 1000000, 229968);
    $display("Test99 completed");
    $display("SUCCESS!");
end
endmodule
